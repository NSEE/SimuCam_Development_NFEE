package rmap_target_read_reply_data_data_pkg is
	
end package rmap_target_read_reply_data_data_pkg;

package body rmap_target_read_reply_data_data_pkg is
	
end package body rmap_target_read_reply_data_data_pkg;
