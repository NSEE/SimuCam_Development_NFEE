// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:51:50 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GwN/QFKroYnPE3m0JowK5DUP6GxDdxd715Y20aE62Q7AlTL4cYVsayTORHVScZUw
ExVSM2EqUeXOoiV8MW96/kgCFckGoqMDYiMKeE0I8Zpk/TSfRQ7yib0C7bgx7hIE
FoEgasG8wk6+Ic8g9AZdcq3Pptt6ArtR+CtWD+p36dM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5344)
Rfaj5Cmj+1Z5UZmU+hb0a56+TfyNqHUZe2jLFuikqw0vi8OhTrj+fPfC7YfrhKMF
At5Ao3ajLNX4f/h4dz47PCQMDmu2akjuLI4P8H+rOQnN1EDCSNYyfWAcHMmTUlwj
IYjq14SkFwcaHZ71GvTciAkUY6Fok//b1pbvQ4a5pdq9eImbUtgq0xh9MEK0fvN6
vwY6If7RaLBACgVyatXIns9Cb7lIi9LPxdoepCWFNK3onPJkGbuWjuHeXOLrjXoH
BHYfNVCkzYNypFBw+TOEquBlxOJlliw+8pgUXwa60ghvqPIHC/55KxWBFz0S7U0z
Uc+2OX5/YFQZp1Jz988MBkOu9ZLUafiEjhP3zAaRaPcMxO/3HprTKPRhGAS1OrGq
0/6HIjlf8HFvGk5OFWH8mQI6R36kQAgGqO13yuVQLLLGK065Uj4dzAOA6z+0WURJ
nlxp9QbdJsbbuqoM1DPg6t61mUCuyLRLmkKDpYX+tgtDgljShCC2lq/hZEOLyTcC
mQ/J09UFcq4ldRVPZS84JP3sZQ2sCHj7Qjb1n2sLocgxvrkRCnu9XcXCPU1Hfe/y
mlkKM5U4bZSEWW8HWPlAGeeY447nhorzvvZXkiPNWTSCS/k02t2+Ou+Nke6yxPcv
nM6T4cMJlNZdpDgFoehxg9bNN4TEx+MupMhlICVjq9/QqeGP39Kg+hJyhZKk3vEF
zptS5AaWU40rWuxNp7kt8rxSLeqPlPD9xZnOHWMc6JUFp9Vw1HuBzOOFxC9Ie3/Z
+iNrDlUxREiB33MP2w2r7QRBnbhqCrpLW/xmMF7bEA6peHkLuGpMxUw05hH0ZmyU
aal8ri2UykYl+H5zRt+ZlioAaME8d7ecFaBTBApudRlCcpDZrT6qBrW6PbYVmB2f
zoIyF8qbIkG+k489YhGvL4162wZnwGP5ssqbj8UC7eEA9kPMM46RnZ8DPQWgT5OT
ygjjMhxbU4NLRifXgQU+8WuPBW8LhQV5UJgVaTvCoKTzx2pBlBTG0pvgTboyN1Xi
S+45wejRgHziuvbQOYoaeDzrnxPVtFGGoGOpDPTPjrEekRiorL4Msa1i8LZskzJR
9Fzc82ZVxAD6FuvXUlVesgpyFHNxCntlhc2q4pE+fe58dD6a+NB9A9ZiA5/J05hU
ejXZHCnGX7D2rymsB1Xzx5gcx0dOIOJcc3rWKOKRP0WC+C9pfHhc98So9hNHHDj1
DqjXL9JbcEs5aD9A+o+Z0MHA1nE20Hr9O6ZeVqZnT7DREcNODo5QcVBAY2Xq8kfC
K7u2WF9vUb097ScHH6iOhs0bA7f4emVfLZA3CJr1Kfmefp4WLA8eDutH4wBA2Jot
gi1BgkvccGDGt/uiozpuWHtIytNd1484l+BQOTLMJTFlvRTiaTltRuGemReBdyIf
WjShLQIOwu++cFdu8GiON1ILeJ0kh8DQcfHw/Do+AEDaiKwu2X3xoWu2t7UloWnR
D/nKR3BznWYYi2lyiZ8YwqsREBBB8gEIQWWiEDB+6W0JqWnHlF9+jES0IjvWSVI6
Qt+AkJ54j0ui6kmhl3Gi5ayq0EoMq55Ztvq6Vpb37j3on7pywozbXC9/tUaCf5NK
Au6ZDPt828fLvrjS17/YEmeOHTck01iLbgWoA0RaojrFlTWbhozc6rTaCthve43C
UfRDqW3Z1YMv94tplN3SfWjGNLjpHanSc4jgKQzJksqzZUkI9NXt9ZwdPX8T1riJ
UcnCkC/LzA0VNg2lnfUJB61Yk2vyY7oGuvq8Tb+1w4WSBPYgPVL7nXmhauPmGVnK
fM8tj+2Md5BGCS0trTjET0ybaCMXD6o4qlYgFjGAS9WEO/LtjRWI9EWAKqhDLBlP
ieWWgIw0G/4WZHxwTmJtJAZbSXUWTF3QFn1yhI2VZLWI1Cwi1015LdXWnLR7KVFk
BAbjQITzEfS2gPQkfGIlTiMzfJiGZNzb2gho12AHvo5XqEKuQxiP6BQmvEnZsy0A
jBqIEnD5MfgPnpWpX8MDonA1osNA+Zgk2qE8B4ugBzhlNZRCJj5GV5I2y0gCN+rh
iqBkCkotzH8gRgc/GkJ2n8sNbai65fy5cFTg3p9V/yZnO0VUeKSjG7yLXGDuOqM0
Oxd3/Xys37uvvEwxVLiNSKjjyCI2hng97bX6gJWBmCumCTzz7MX+z3ZkO6fKsya+
qdnd+pSCth8DjOu+toBhQBTb7379475OEYKOKSevWLOdV7ZIHgpRcZLqyqxEXwk8
gLzRPUbBVb6Q6RRVEx7/YR2hjSCacT36CE/A/mnrkOEAUvnZJ4zNRzPc7MndaKUj
10h+LavfKS9BQ2itsBe7dPUmV5ogCW4WuQ5+KBbGXkKSu8IZXTVbCRrIsqWJnxCd
RJ5diLtREmpJFpqDosGrpakDx0DznGF6IpkFlWaL56xQLDA35Dn+wmdm+Kwt3E7Y
P305GRPULKGZOWOThm7rNIIyxuSg0DoA80zisRzcpxS4GaNHN9mSOespw8zHdgSD
DDxcCp1KrsT5KDzzHLWXCXHv/QqQPmpqysx5Cqei/JGIhBETd5Zed/Td7Dx1buiF
aNkONEmEp6ec6XnHP1AastPI7vdBHe3BDF+4fBF/+zmEr6g86VgHVZkSRR130UjD
yxbT6KC0u1c++psuonmXtV5G2WODQdHAO9+W4rEYhrqm7QCK7k6/LJgtb8VLQFWB
tp8WUeGtt3AtUX0yY0lfUOhAik99nqFkR4SysoE7JNuJcAJ3geuJ0m6+6iUYIAVD
/UNJIROZNkslXkypF57zwboq8/EbFGVsTfDzr7fu8hLapfMXEUAocbwqO4mTJ248
jgEDeCF386dxugao0zP0TImTf4QI3pvmcLFCOLXDsGBVF3COtojQmtEK2EXgCbpj
Bnmk/CoJ3VXC9wzKPgaVXbOdQFZE+fgFs/eJhbKNO/3rlQhJlRdpohQAYbuK04tm
w8z4h5QwTOg/lzf897C6gYsrrIgELhJivZ4RQz+z1s3FWAFSI7Kl3RffXML72bEg
b5qxzB77qNCPBGfFpQv2WHZ4GctBp2VhzXxp/LfZBUqYAq34RIFBe7cDtK8V+ukh
ahfJ0b08MTFLtWoKFQxvxHIgms15pcCW4cG6urJCjp2k+wkTGT2X6FemKKVyeavK
k9KgkJpt8q2FsLcRuxDdPIPx56RX6mFyVCc8klnEno6QVpfkL92wt133WWdGQTnJ
NZsf6YVIDpSKn+sxlPDnscAc+ezun/WIgjR1uCnQ+Tfq8LlLDyD5UQHU0qJ8s//k
cG2NttF7qedrpPhutqJzFhW0ihYFxQmEpfHdaiHXCKTov58eyy3NQKV562WYrw91
3EBn9RWBj+wcFlbg5qU4nWYSB4qgOQ71q8SvsLU/IvsJ2um1xYqS4cgXXOpXneuH
ilYw92tMO7ybXo8OxIzZPHlnaGSwMR8KIUeniM5LhyNc0fLJ4rDlnzzzb5MopDzB
KA1P9XPXs8XjnWtwH4p8V+zTN0cQm65+9+j3cw0P1LA4TDngCCRJLspYLecxsouT
D0PR6weIiV3aQvK8J8lumA6hFtJ6HMHONFqIH0tClSf+pQaHkJMEIWFJ4W+JF63G
q6VvJy1sRPTl6d2KCufSu1jJkK9qSfiWDYNVsq4ZrXZ7PbixlkbiwFjfH0toljyg
wa8qdKDQ7Z/bB/O+ut9WNhc/etnzSOXyFLrmJfTpAjhCT8qeWCgqhsTudoEHm3Oe
E2iM9VjP8K7pNgCupmoJ00BcF11zPc76fxO1kRWqVfj5KM3aqtZNICc6PnHGwMkI
ybLRFLJdHy/GsTFoS79OeCuHNwflQHVinpqc05X2wVeRTRakalxNmotYlnqysG1C
4GreHR5rYVHIv7QH5HhP084JIRFf2yZtVJQbkYJ27sgHbXG5m6XBF/tQqi/kQG8Q
QnaOFIdRxozAnkaDNKXJ/rofHaFJ+Q9lGIjocb2AkWs9+k3MZhaEBBq7bSpCCFRg
alait8NO91b9rLmlolzsAyLTtdYwFhVyPp2KrQRkVKQJ50gTpdW/RsrePJJ/lpnA
CH2frmqbsbDGakZOnRh7zdkQYOaGTbtwcLk2cMytLkb9MmzARj3D/sc4S0pwe/HD
oyfFVl1zvZkH9kp75/MUV63tcg5D6TRKt/y631+jCSuIp1aLZInHQSIyYsraQ4fv
BNemjtDuR1ohJEJMjrGXHU0QAdIxMmN7xsi0xQ3Sdzs4zxD/ncbNAd/M0YJY6SQ7
uZzXvVBv75LejBq7WA77ouXK0CuRu6CEC8UOqgTpEZN0mlNVCDQcRGxXXfTrBxIV
K4nf4F2eixDhAgeqzHN2Z0GsWIC57W1dXS8VRHwtLF8u+QhDope+VWcyrrTRMimQ
6ka04XX+THBVRezOED1zeKo3AEXZnL/Ihu92mMh69L6jK1U+2SHswEOb5U49e8K5
uVmtX9367/hk99pq9vJWbJNwdrTEyeS1Xs1vl1LmpLcBBKsOUA6BLziX/gwgh9r6
i+rTT0l7sSCBM1JR8qVEpuSdoWfTkm9I/mvPsaARcNZRnC29vKNuAH7k4KRsAv8Y
fMIKy8p5Aukk/agk1J/Ux+F2LRkQiPQJRPCV28kK6iYm+ufqAmkN/yNv8e6yX03C
69KAgIwHL/jHM24JAb9h3/uwLXscs0w63jJGhBp1IMx/DMbIoPOX8owSRzcIxMx8
DYw1pf1g2PY3j4aVZBcdWwP1FuPwIfrJO5+9wayOw/jH02oRu7FRoMTcfPx/vQTz
bMaalVixm1Rk1zXwJLXJZyGzai4NNVeUNbYrGjI7f2cZy9/rKg6ADG6b+8SAWYGR
BTmxJMfOAErDZmIde0BW9mIEb+9cUXaZO9blnUj4qN9wrQeIWy/VphHTn1sgJQDk
DqW4prTz/wjTvGxDGlqd7p19O5q+uR5bcxSV69DDBy8ZK4XafoPgq9P0RMUBEmai
5BHXvucryNzPPNykMiaFrlmLdd4pLzBnQ49OK5zV2OuUOvUFnb30g+Hj9tI+hX+c
zJp/9KoEjjED242Fp5OF90ixWnXLBhsU05YfstyXohppGnzKT5hvDYwiJlyP0Le+
DHzLQW6ZZJI0gg2xdQ4RgCZbDFeeefvetXb+BzM0reFDaZpfN2ZLtQPCuNVJ+imL
gcC4xyJQ9ax0ZPoL2x9oU3gbHdLRXODy0TEEuxt9+CoH0NIDYVhf+stYBEAju9AC
1Fma0ZACZ7Y9vV3NQak26+NeHZKpUegki0c4p1cBRLJqRb0M+EAywZbrETZ37Vam
0xLEEU1jpHPtzagEiQxIhoAcwHGPvNYOTLWr9afCJNybyxg1K3nPXk6StFaxuJeL
N5OPdkdoF8QnTDWQ0Yngpfyl+rh/JXczRNUy4ZKeP1LQ9ePapbp2XlUHgYWtZN4E
lh2a9KLQDFf8h5Ius8EyE218dSg7S4fOJVs1bUrLkpczt+doyBrmdpYJGK7K9+jl
H19OfrzBRUvIL+G605Ys0VwBN0J9NR/y3QoAfUisWkQi3bVn8VuglHztxRb0m5uH
cRhlrYE6WWoUqlVG79tUjSsKpHQZOLDKxRuqgo/eFtWGO9QZhQjNV8zVb2/R2yhg
N+Lkb3Qm5dEZoui9WS8NhMnK9cG5xOz4LpY/2LVO2nYlQ6reOwxQeM5Tdo8JUHrF
UnxT8F+KBdsv1Td+nHz2A5YCELQQK3BN41r/M6EjagTG3JGvZjeCyk1rmB884/Kx
IhYusrO954LC+Pp70wMLTY+AmMk3s61E6kY4fyGotg2nLGXAe0y6zKSP96BZT+Hw
RlHoRRr55y3hSEYocMwb2LUqTLmBIssaWupxrdKEH1hEOLI+4LbzqRC+RmKtLnFb
Ub5+jylgSuumP4wyes4nvT1eHuR+tr37wTaQ8DosL0ajJM2LyPavyq7Kb43RRH+T
/UuvG0rtBhTymeG54k8RwFHEAwgEFMsKm5V00nawmjK39JGUQLNQC5bColsOw8R/
VZZHj7cSh6tjC33rBeKo1HDzofFZoDyaSq//57+b989/2vUmz6839jvCHncr0WhL
5Os0hjRJ2giRK4ktgyy2Cf3Ir5O7mXzEhXXMtlaGRYJkuf1Lqb3smGF4vNkh5uVa
RBGAZl2wlTnijUxgmSFw2GT5HrliaVxepGz4OA3uG0/T5CKgxBvqiNCFgS8ZX7Eb
+1dOauwLGIbIwm/kULRl3GA1wUE7Bi1+HzYrdz8NEdNpy9mQv8JxOxWBGzx7+Kc9
hL6xkA4eC9Ayz/nxv7Wu2iWeLzKH1+5UA1zQ2yyQD7kM1tmOIEaciwyBhNvpAwQn
zlSA7Qm3kJpgemHwi4UDo1D2pR6Pp6VcK80LuK0UIGqC8IdAMW7qCOG27QyFuMRe
PFrU8Q0d2GdIayGmpUvRK4I2/O02fHG7K6Pga3uuO0ApqKtvITxnmczSjv1NFokg
zBfq9nMlszElByamiXoANEkTaWbHJTds13+P9KkKIe0qCYjv3ZRxHr9pVzNq+b4c
O3yzcwObLVYRtugArI0ejE0SxOhaHQkWsVl9wePASL9+/DP0LyNV+K+b7WOp5GSl
VJvuWvhnqXKAW2wNzLNFM3zstE+tFUou6DebmLXgT2maOeFZJZ9xB9FQq76nSscQ
p7VNHcIdXL1HMedulpYwEw8nUH1lrFUqi+oxSAPWFfRBAXPgzV82SWrETa3OqfuH
nPBOBGGcubYieB6JSZMHaLQ32JSZolzzFzfDlSamhJF0aFfq+5GA1DYjQ6hT0jSy
jEh6w/NLhH0THN+eb0IMh9/5lkrCcp2l2+dykMyyd9gDiBdpDkYqCxPGv/7mAlc/
fOVhvhmqJBegbsBHlfJi3rX+l1qvJkJxD+IyxZ1JQbs8RxUPILz0YG/pAzxm53pP
fbS1MsQklVpTWmbEq8thYb/fRdiyUVmIxmyCRK3uqzZeObHNnp1lor4+cbyx9EgO
UnUEryZ+peL/zqV0LTIXskR4vBKYVDqz5pk8LJoVMQwOz6II528b6swdP+GaJlb8
1IdK/ZSXp7kyW4s6EilwBZKYb3zZaAfJvy0nNyUeKdIXP5mEYG30ywWnv0inH0gw
hDOcKxSbsvA0gEXyMuVUf4NSgP7nK+bQ6pJd5Lhy0Ev3BcxNFwBIYe2x40Cb4VgI
x3mpmWD0jwr63OWQVxHDbw==
`pragma protect end_protected
