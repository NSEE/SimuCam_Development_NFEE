// MebX_Qsys_Project.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module MebX_Qsys_Project (
		input  wire [3:0]  button_export,                                               //                               button.export
		input  wire        clk50_clk,                                                   //                                clk50.clk
		output wire [7:0]  comm_a_measurements_conduit_end_measurements_channel_signal, //      comm_a_measurements_conduit_end.measurements_channel_signal
		input  wire        comm_a_sync_end_sync_channel_signal,                         //                      comm_a_sync_end.sync_channel_signal
		output wire [7:0]  comm_b_measurements_conduit_end_measurements_channel_signal, //      comm_b_measurements_conduit_end.measurements_channel_signal
		input  wire        comm_b_sync_end_sync_channel_signal,                         //                      comm_b_sync_end.sync_channel_signal
		output wire [7:0]  comm_c_measurements_conduit_end_measurements_channel_signal, //      comm_c_measurements_conduit_end.measurements_channel_signal
		input  wire        comm_c_sync_end_sync_channel_signal,                         //                      comm_c_sync_end.sync_channel_signal
		output wire [7:0]  comm_d_measurements_conduit_end_measurements_channel_signal, //      comm_d_measurements_conduit_end.measurements_channel_signal
		input  wire        comm_d_sync_end_sync_channel_signal,                         //                      comm_d_sync_end.sync_channel_signal
		output wire [7:0]  comm_e_measurements_conduit_end_measurements_channel_signal, //      comm_e_measurements_conduit_end.measurements_channel_signal
		input  wire        comm_e_sync_end_sync_channel_signal,                         //                      comm_e_sync_end.sync_channel_signal
		output wire [7:0]  comm_f_measurements_conduit_end_measurements_channel_signal, //      comm_f_measurements_conduit_end.measurements_channel_signal
		input  wire        comm_f_sync_end_sync_channel_signal,                         //                      comm_f_sync_end.sync_channel_signal
		output wire        csense_adc_fo_export,                                        //                        csense_adc_fo.export
		output wire [1:0]  csense_cs_n_export,                                          //                          csense_cs_n.export
		output wire        csense_sck_export,                                           //                           csense_sck.export
		output wire        csense_sdi_export,                                           //                           csense_sdi.export
		input  wire        csense_sdo_export,                                           //                           csense_sdo.export
		output wire [3:0]  ctrl_io_lvds_export,                                         //                         ctrl_io_lvds.export
		input  wire [7:0]  dip_export,                                                  //                                  dip.export
		input  wire        ext_export,                                                  //                                  ext.export
		input  wire        ftdi_clk_clk,                                                //                             ftdi_clk.clk
		output wire [7:0]  led_de4_export,                                              //                              led_de4.export
		output wire [20:0] led_painel_export,                                           //                           led_painel.export
		output wire        m1_ddr2_i2c_scl_export,                                      //                      m1_ddr2_i2c_scl.export
		inout  wire        m1_ddr2_i2c_sda_export,                                      //                      m1_ddr2_i2c_sda.export
		output wire [13:0] m1_ddr2_memory_mem_a,                                        //                       m1_ddr2_memory.mem_a
		output wire [2:0]  m1_ddr2_memory_mem_ba,                                       //                                     .mem_ba
		output wire [1:0]  m1_ddr2_memory_mem_ck,                                       //                                     .mem_ck
		output wire [1:0]  m1_ddr2_memory_mem_ck_n,                                     //                                     .mem_ck_n
		output wire [1:0]  m1_ddr2_memory_mem_cke,                                      //                                     .mem_cke
		output wire [1:0]  m1_ddr2_memory_mem_cs_n,                                     //                                     .mem_cs_n
		output wire [7:0]  m1_ddr2_memory_mem_dm,                                       //                                     .mem_dm
		output wire [0:0]  m1_ddr2_memory_mem_ras_n,                                    //                                     .mem_ras_n
		output wire [0:0]  m1_ddr2_memory_mem_cas_n,                                    //                                     .mem_cas_n
		output wire [0:0]  m1_ddr2_memory_mem_we_n,                                     //                                     .mem_we_n
		inout  wire [63:0] m1_ddr2_memory_mem_dq,                                       //                                     .mem_dq
		inout  wire [7:0]  m1_ddr2_memory_mem_dqs,                                      //                                     .mem_dqs
		inout  wire [7:0]  m1_ddr2_memory_mem_dqs_n,                                    //                                     .mem_dqs_n
		output wire [1:0]  m1_ddr2_memory_mem_odt,                                      //                                     .mem_odt
		input  wire        m1_ddr2_memory_pll_ref_clk_clk,                              //           m1_ddr2_memory_pll_ref_clk.clk
		output wire        m1_ddr2_memory_status_local_init_done,                       //                m1_ddr2_memory_status.local_init_done
		output wire        m1_ddr2_memory_status_local_cal_success,                     //                                     .local_cal_success
		output wire        m1_ddr2_memory_status_local_cal_fail,                        //                                     .local_cal_fail
		input  wire        m1_ddr2_oct_rdn,                                             //                          m1_ddr2_oct.rdn
		input  wire        m1_ddr2_oct_rup,                                             //                                     .rup
		output wire        m2_ddr2_i2c_scl_export,                                      //                      m2_ddr2_i2c_scl.export
		inout  wire        m2_ddr2_i2c_sda_export,                                      //                      m2_ddr2_i2c_sda.export
		output wire [13:0] m2_ddr2_memory_mem_a,                                        //                       m2_ddr2_memory.mem_a
		output wire [2:0]  m2_ddr2_memory_mem_ba,                                       //                                     .mem_ba
		output wire [1:0]  m2_ddr2_memory_mem_ck,                                       //                                     .mem_ck
		output wire [1:0]  m2_ddr2_memory_mem_ck_n,                                     //                                     .mem_ck_n
		output wire [1:0]  m2_ddr2_memory_mem_cke,                                      //                                     .mem_cke
		output wire [1:0]  m2_ddr2_memory_mem_cs_n,                                     //                                     .mem_cs_n
		output wire [7:0]  m2_ddr2_memory_mem_dm,                                       //                                     .mem_dm
		output wire [0:0]  m2_ddr2_memory_mem_ras_n,                                    //                                     .mem_ras_n
		output wire [0:0]  m2_ddr2_memory_mem_cas_n,                                    //                                     .mem_cas_n
		output wire [0:0]  m2_ddr2_memory_mem_we_n,                                     //                                     .mem_we_n
		inout  wire [63:0] m2_ddr2_memory_mem_dq,                                       //                                     .mem_dq
		inout  wire [7:0]  m2_ddr2_memory_mem_dqs,                                      //                                     .mem_dqs
		inout  wire [7:0]  m2_ddr2_memory_mem_dqs_n,                                    //                                     .mem_dqs_n
		output wire [1:0]  m2_ddr2_memory_mem_odt,                                      //                                     .mem_odt
		input  wire        m2_ddr2_memory_dll_sharing_dll_pll_locked,                   //           m2_ddr2_memory_dll_sharing.dll_pll_locked
		output wire [5:0]  m2_ddr2_memory_dll_sharing_dll_delayctrl,                    //                                     .dll_delayctrl
		output wire        m2_ddr2_memory_pll_sharing_pll_mem_clk,                      //           m2_ddr2_memory_pll_sharing.pll_mem_clk
		output wire        m2_ddr2_memory_pll_sharing_pll_write_clk,                    //                                     .pll_write_clk
		output wire        m2_ddr2_memory_pll_sharing_pll_locked,                       //                                     .pll_locked
		output wire        m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk,        //                                     .pll_write_clk_pre_phy_clk
		output wire        m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk,                 //                                     .pll_addr_cmd_clk
		output wire        m2_ddr2_memory_pll_sharing_pll_avl_clk,                      //                                     .pll_avl_clk
		output wire        m2_ddr2_memory_pll_sharing_pll_config_clk,                   //                                     .pll_config_clk
		output wire        m2_ddr2_memory_status_local_init_done,                       //                m2_ddr2_memory_status.local_init_done
		output wire        m2_ddr2_memory_status_local_cal_success,                     //                                     .local_cal_success
		output wire        m2_ddr2_memory_status_local_cal_fail,                        //                                     .local_cal_fail
		input  wire        m2_ddr2_oct_rdn,                                             //                          m2_ddr2_oct.rdn
		input  wire        m2_ddr2_oct_rup,                                             //                                     .rup
		input  wire        rs232_uart_rxd,                                              //                           rs232_uart.rxd
		output wire        rs232_uart_txd,                                              //                                     .txd
		input  wire        rst_reset_n,                                                 //                                  rst.reset_n
		input  wire        rst_controller_conduit_reset_input_t_reset_input_signal,     //   rst_controller_conduit_reset_input.t_reset_input_signal
		output wire        rst_controller_conduit_simucam_reset_t_simucam_reset_signal, // rst_controller_conduit_simucam_reset.t_simucam_reset_signal
		input  wire        rtcc_alarm_export,                                           //                           rtcc_alarm.export
		output wire        rtcc_cs_n_export,                                            //                            rtcc_cs_n.export
		output wire        rtcc_sck_export,                                             //                             rtcc_sck.export
		output wire        rtcc_sdi_export,                                             //                             rtcc_sdi.export
		input  wire        rtcc_sdo_export,                                             //                             rtcc_sdo.export
		inout  wire        sd_card_ip_b_SD_cmd,                                         //                           sd_card_ip.b_SD_cmd
		inout  wire        sd_card_ip_b_SD_dat,                                         //                                     .b_SD_dat
		inout  wire        sd_card_ip_b_SD_dat3,                                        //                                     .b_SD_dat3
		output wire        sd_card_ip_o_SD_clock,                                       //                                     .o_SD_clock
		input  wire        sd_card_wp_n_io_export,                                      //                      sd_card_wp_n_io.export
		input  wire        spwc_a_enable_spw_rx_enable_signal,                          //                        spwc_a_enable.spw_rx_enable_signal
		input  wire        spwc_a_enable_spw_tx_enable_signal,                          //                                     .spw_tx_enable_signal
		output wire        spwc_a_leds_spw_red_status_led_signal,                       //                          spwc_a_leds.spw_red_status_led_signal
		output wire        spwc_a_leds_spw_green_status_led_signal,                     //                                     .spw_green_status_led_signal
		input  wire        spwc_a_lvds_spw_lvds_data_in_signal,                         //                          spwc_a_lvds.spw_lvds_data_in_signal
		output wire        spwc_a_lvds_spw_lvds_data_out_signal,                        //                                     .spw_lvds_data_out_signal
		output wire        spwc_a_lvds_spw_lvds_strobe_out_signal,                      //                                     .spw_lvds_strobe_out_signal
		input  wire        spwc_a_lvds_spw_lvds_strobe_in_signal,                       //                                     .spw_lvds_strobe_in_signal
		input  wire        spwc_b_enable_spw_rx_enable_signal,                          //                        spwc_b_enable.spw_rx_enable_signal
		input  wire        spwc_b_enable_spw_tx_enable_signal,                          //                                     .spw_tx_enable_signal
		output wire        spwc_b_leds_spw_red_status_led_signal,                       //                          spwc_b_leds.spw_red_status_led_signal
		output wire        spwc_b_leds_spw_green_status_led_signal,                     //                                     .spw_green_status_led_signal
		input  wire        spwc_b_lvds_spw_lvds_data_in_signal,                         //                          spwc_b_lvds.spw_lvds_data_in_signal
		output wire        spwc_b_lvds_spw_lvds_data_out_signal,                        //                                     .spw_lvds_data_out_signal
		output wire        spwc_b_lvds_spw_lvds_strobe_out_signal,                      //                                     .spw_lvds_strobe_out_signal
		input  wire        spwc_b_lvds_spw_lvds_strobe_in_signal,                       //                                     .spw_lvds_strobe_in_signal
		input  wire        spwc_c_enable_spw_rx_enable_signal,                          //                        spwc_c_enable.spw_rx_enable_signal
		input  wire        spwc_c_enable_spw_tx_enable_signal,                          //                                     .spw_tx_enable_signal
		output wire        spwc_c_leds_spw_red_status_led_signal,                       //                          spwc_c_leds.spw_red_status_led_signal
		output wire        spwc_c_leds_spw_green_status_led_signal,                     //                                     .spw_green_status_led_signal
		input  wire        spwc_c_lvds_spw_lvds_data_in_signal,                         //                          spwc_c_lvds.spw_lvds_data_in_signal
		output wire        spwc_c_lvds_spw_lvds_data_out_signal,                        //                                     .spw_lvds_data_out_signal
		output wire        spwc_c_lvds_spw_lvds_strobe_out_signal,                      //                                     .spw_lvds_strobe_out_signal
		input  wire        spwc_c_lvds_spw_lvds_strobe_in_signal,                       //                                     .spw_lvds_strobe_in_signal
		input  wire        spwc_d_enable_spw_rx_enable_signal,                          //                        spwc_d_enable.spw_rx_enable_signal
		input  wire        spwc_d_enable_spw_tx_enable_signal,                          //                                     .spw_tx_enable_signal
		output wire        spwc_d_leds_spw_red_status_led_signal,                       //                          spwc_d_leds.spw_red_status_led_signal
		output wire        spwc_d_leds_spw_green_status_led_signal,                     //                                     .spw_green_status_led_signal
		input  wire        spwc_d_lvds_spw_lvds_data_in_signal,                         //                          spwc_d_lvds.spw_lvds_data_in_signal
		output wire        spwc_d_lvds_spw_lvds_data_out_signal,                        //                                     .spw_lvds_data_out_signal
		output wire        spwc_d_lvds_spw_lvds_strobe_out_signal,                      //                                     .spw_lvds_strobe_out_signal
		input  wire        spwc_d_lvds_spw_lvds_strobe_in_signal,                       //                                     .spw_lvds_strobe_in_signal
		input  wire        spwc_e_enable_spw_rx_enable_signal,                          //                        spwc_e_enable.spw_rx_enable_signal
		input  wire        spwc_e_enable_spw_tx_enable_signal,                          //                                     .spw_tx_enable_signal
		output wire        spwc_e_leds_spw_red_status_led_signal,                       //                          spwc_e_leds.spw_red_status_led_signal
		output wire        spwc_e_leds_spw_green_status_led_signal,                     //                                     .spw_green_status_led_signal
		input  wire        spwc_e_lvds_spw_lvds_data_in_signal,                         //                          spwc_e_lvds.spw_lvds_data_in_signal
		output wire        spwc_e_lvds_spw_lvds_data_out_signal,                        //                                     .spw_lvds_data_out_signal
		output wire        spwc_e_lvds_spw_lvds_strobe_out_signal,                      //                                     .spw_lvds_strobe_out_signal
		input  wire        spwc_e_lvds_spw_lvds_strobe_in_signal,                       //                                     .spw_lvds_strobe_in_signal
		input  wire        spwc_f_enable_spw_rx_enable_signal,                          //                        spwc_f_enable.spw_rx_enable_signal
		input  wire        spwc_f_enable_spw_tx_enable_signal,                          //                                     .spw_tx_enable_signal
		output wire        spwc_f_leds_spw_red_status_led_signal,                       //                          spwc_f_leds.spw_red_status_led_signal
		output wire        spwc_f_leds_spw_green_status_led_signal,                     //                                     .spw_green_status_led_signal
		input  wire        spwc_f_lvds_spw_lvds_data_in_signal,                         //                          spwc_f_lvds.spw_lvds_data_in_signal
		output wire        spwc_f_lvds_spw_lvds_data_out_signal,                        //                                     .spw_lvds_data_out_signal
		output wire        spwc_f_lvds_spw_lvds_strobe_out_signal,                      //                                     .spw_lvds_strobe_out_signal
		input  wire        spwc_f_lvds_spw_lvds_strobe_in_signal,                       //                                     .spw_lvds_strobe_in_signal
		input  wire        spwc_g_enable_spw_rx_enable_signal,                          //                        spwc_g_enable.spw_rx_enable_signal
		input  wire        spwc_g_enable_spw_tx_enable_signal,                          //                                     .spw_tx_enable_signal
		output wire        spwc_g_leds_spw_red_status_led_signal,                       //                          spwc_g_leds.spw_red_status_led_signal
		output wire        spwc_g_leds_spw_green_status_led_signal,                     //                                     .spw_green_status_led_signal
		input  wire        spwc_g_lvds_spw_lvds_data_in_signal,                         //                          spwc_g_lvds.spw_lvds_data_in_signal
		output wire        spwc_g_lvds_spw_lvds_data_out_signal,                        //                                     .spw_lvds_data_out_signal
		output wire        spwc_g_lvds_spw_lvds_strobe_out_signal,                      //                                     .spw_lvds_strobe_out_signal
		input  wire        spwc_g_lvds_spw_lvds_strobe_in_signal,                       //                                     .spw_lvds_strobe_in_signal
		input  wire        spwc_h_enable_spw_rx_enable_signal,                          //                        spwc_h_enable.spw_rx_enable_signal
		input  wire        spwc_h_enable_spw_tx_enable_signal,                          //                                     .spw_tx_enable_signal
		output wire        spwc_h_leds_spw_red_status_led_signal,                       //                          spwc_h_leds.spw_red_status_led_signal
		output wire        spwc_h_leds_spw_green_status_led_signal,                     //                                     .spw_green_status_led_signal
		input  wire        spwc_h_lvds_spw_lvds_data_in_signal,                         //                          spwc_h_lvds.spw_lvds_data_in_signal
		output wire        spwc_h_lvds_spw_lvds_data_out_signal,                        //                                     .spw_lvds_data_out_signal
		output wire        spwc_h_lvds_spw_lvds_strobe_out_signal,                      //                                     .spw_lvds_strobe_out_signal
		input  wire        spwc_h_lvds_spw_lvds_strobe_in_signal,                       //                                     .spw_lvds_strobe_in_signal
		input  wire        sync_in_conduit,                                             //                              sync_in.conduit
		output wire        sync_out_conduit,                                            //                             sync_out.conduit
		output wire        sync_spw1_conduit,                                           //                            sync_spw1.conduit
		output wire        sync_spw2_conduit,                                           //                            sync_spw2.conduit
		output wire        sync_spw3_conduit,                                           //                            sync_spw3.conduit
		output wire        sync_spw4_conduit,                                           //                            sync_spw4.conduit
		output wire        sync_spw5_conduit,                                           //                            sync_spw5.conduit
		output wire        sync_spw6_conduit,                                           //                            sync_spw6.conduit
		output wire        sync_spw7_conduit,                                           //                            sync_spw7.conduit
		output wire        sync_spw8_conduit,                                           //                            sync_spw8.conduit
		output wire        temp_scl_export,                                             //                             temp_scl.export
		inout  wire        temp_sda_export,                                             //                             temp_sda.export
		output wire        timer_1ms_external_port_export,                              //              timer_1ms_external_port.export
		output wire        timer_1us_external_port_export,                              //              timer_1us_external_port.export
		output wire [25:0] tristate_conduit_tcm_address_out,                            //                     tristate_conduit.tcm_address_out
		output wire [0:0]  tristate_conduit_tcm_read_n_out,                             //                                     .tcm_read_n_out
		output wire [0:0]  tristate_conduit_tcm_write_n_out,                            //                                     .tcm_write_n_out
		inout  wire [15:0] tristate_conduit_tcm_data_out,                               //                                     .tcm_data_out
		output wire [0:0]  tristate_conduit_tcm_chipselect_n_out,                       //                                     .tcm_chipselect_n_out
		inout  wire [31:0] umft601a_pins_umft_data_signal,                              //                        umft601a_pins.umft_data_signal
		output wire        umft601a_pins_umft_reset_n_signal,                           //                                     .umft_reset_n_signal
		input  wire        umft601a_pins_umft_rxf_n_signal,                             //                                     .umft_rxf_n_signal
		input  wire        umft601a_pins_umft_clock_signal,                             //                                     .umft_clock_signal
		inout  wire        umft601a_pins_umft_wakeup_n_signal,                          //                                     .umft_wakeup_n_signal
		inout  wire [3:0]  umft601a_pins_umft_be_signal,                                //                                     .umft_be_signal
		input  wire        umft601a_pins_umft_txe_n_signal,                             //                                     .umft_txe_n_signal
		inout  wire [1:0]  umft601a_pins_umft_gpio_bus_signal,                          //                                     .umft_gpio_bus_signal
		output wire        umft601a_pins_umft_wr_n_signal,                              //                                     .umft_wr_n_signal
		output wire        umft601a_pins_umft_rd_n_signal,                              //                                     .umft_rd_n_signal
		output wire        umft601a_pins_umft_oe_n_signal,                              //                                     .umft_oe_n_signal
		output wire        umft601a_pins_umft_siwu_n_signal                             //                                     .umft_siwu_n_signal
	);

	wire          m2_ddr2_memory_afi_clk_clk;                                                                // m2_ddr2_memory:afi_clk -> [COMM_Pedreiro_v1_01_1:clock_sink_200_clk, COMM_Pedreiro_v1_01_2:clock_sink_200_clk, COMM_Pedreiro_v1_01_3:clock_sink_200_clk, COMM_Pedreiro_v1_01_4:clock_sink_200_clk, COMM_Pedreiro_v1_01_5:clock_sink_200_clk, COMM_Pedreiro_v1_01_6:clock_sink_200_clk, SpaceWire_Channel_A:clk_200_i, SpaceWire_Channel_B:clk_200_i, SpaceWire_Channel_C:clk_200_i, SpaceWire_Channel_D:clk_200_i, SpaceWire_Channel_E:clk_200_i, SpaceWire_Channel_F:clk_200_i, SpaceWire_Channel_G:clk_200_i, SpaceWire_Channel_H:clk_200_i, mm_interconnect_0:m2_ddr2_memory_afi_clk_clk, rst_controller_010:clk, rst_controller_011:clk, rst_controller_012:clk, rst_controller_013:clk, rst_controller_014:clk, rst_controller_015:clk, rst_controller_016:clk, rst_controller_017:clk, rst_controller_025:clk]
	wire          m2_ddr2_memory_afi_half_clk_clk;                                                           // m2_ddr2_memory:afi_half_clk -> [COMM_Pedreiro_v1_01_1:clock_sink_100_clk, COMM_Pedreiro_v1_01_2:clock_sink_100_clk, COMM_Pedreiro_v1_01_3:clock_sink_100_clk, COMM_Pedreiro_v1_01_4:clock_sink_100_clk, COMM_Pedreiro_v1_01_5:clock_sink_100_clk, COMM_Pedreiro_v1_01_6:clock_sink_100_clk, FTDI_USB3_0:clock_sink_clk, RMAP_Echoing_0:clk_100_i, SpaceWire_Channel_A:clk_100_i, SpaceWire_Channel_B:clk_100_i, SpaceWire_Channel_C:clk_100_i, SpaceWire_Channel_D:clk_100_i, SpaceWire_Channel_E:clk_100_i, SpaceWire_Channel_F:clk_100_i, SpaceWire_Channel_G:clk_100_i, SpaceWire_Channel_H:clk_100_i, SpaceWire_Glutton_0:clk_100_i, clock_bridge_afi_50:s0_clk, ddr2_address_span_extender:clk, ext_flash:clk_clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, irq_synchronizer_004:sender_clk, jtag_uart_0:clk, m1_clock_bridge:s0_clk, mm_interconnect_0:clk_100_clk_clk, mm_interconnect_0:m2_ddr2_memory_afi_half_clk_clk, mm_interconnect_1:clk_100_clk_clk, nios2_gen2_0:clk, onchip_memory:clk, rmap_mem_nfee_comm_1:clk_100_i, rmap_mem_nfee_comm_2:clk_100_i, rmap_mem_nfee_comm_3:clk_100_i, rmap_mem_nfee_comm_4:clk_100_i, rmap_mem_nfee_comm_5:clk_100_i, rmap_mem_nfee_comm_6:clk_100_i, rst_controller_002:clk, rst_controller_003:clk, rst_controller_004:clk, rst_controller_005:clk, rst_controller_006:clk, rst_controller_007:clk, rst_controller_008:clk, rst_controller_009:clk, rst_controller_018:clk, rst_controller_020:clk, rst_controller_022:clk, sysid_qsys:clock, tristate_conduit_bridge_0:clk]
	wire          m1_ddr2_memory_afi_half_clk_clk;                                                           // m1_ddr2_memory:afi_half_clk -> [m1_clock_bridge:m0_clk, mm_interconnect_3:m1_ddr2_memory_afi_half_clk_clk, rst_controller_021:clk]
	wire          comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_e_side_buffer_full_signal;            // COMM_Pedreiro_v1_01_1:channel_hk_err_e_side_buffer_full_o -> rmap_mem_nfee_comm_1:channel_hk_err_e_side_buffer_full_i
	wire          comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_escape_err_signal;               // COMM_Pedreiro_v1_01_1:channel_hk_spw_link_escape_err_o -> rmap_mem_nfee_comm_1:channel_hk_spw_link_escape_err_i
	wire          comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_rmap_target_indicate_signal;              // COMM_Pedreiro_v1_01_1:channel_hk_rmap_target_indicate_o -> rmap_mem_nfee_comm_1:channel_hk_rmap_target_indicate_i
	wire          comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal;             // COMM_Pedreiro_v1_01_1:channel_hk_err_win_wrong_y_coord_o -> rmap_mem_nfee_comm_1:channel_hk_err_win_wrong_y_coord_i
	wire          comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_running_signal;                  // COMM_Pedreiro_v1_01_1:channel_hk_spw_link_running_o -> rmap_mem_nfee_comm_1:channel_hk_spw_link_running_i
	wire          comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_credit_err_signal;               // COMM_Pedreiro_v1_01_1:channel_hk_spw_link_credit_err_o -> rmap_mem_nfee_comm_1:channel_hk_spw_link_credit_err_i
	wire          comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal;             // COMM_Pedreiro_v1_01_1:channel_hk_err_win_wrong_x_coord_o -> rmap_mem_nfee_comm_1:channel_hk_err_win_wrong_x_coord_i
	wire    [7:0] comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_rmap_target_status_signal;                // COMM_Pedreiro_v1_01_1:channel_hk_rmap_target_status_o -> rmap_mem_nfee_comm_1:channel_hk_rmap_target_status_i
	wire          comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_f_side_buffer_full_signal;            // COMM_Pedreiro_v1_01_1:channel_hk_err_f_side_buffer_full_o -> rmap_mem_nfee_comm_1:channel_hk_err_f_side_buffer_full_i
	wire    [5:0] comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_timecode_time_signal;                     // COMM_Pedreiro_v1_01_1:channel_hk_timecode_time_o -> rmap_mem_nfee_comm_1:channel_hk_timecode_time_i
	wire          comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_parity_err_signal;               // COMM_Pedreiro_v1_01_1:channel_hk_spw_link_parity_err_o -> rmap_mem_nfee_comm_1:channel_hk_spw_link_parity_err_i
	wire          comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_disconnect_signal;               // COMM_Pedreiro_v1_01_1:channel_hk_spw_link_disconnect_o -> rmap_mem_nfee_comm_1:channel_hk_spw_link_disconnect_i
	wire          comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal;              // COMM_Pedreiro_v1_01_1:channel_hk_err_invalid_ccd_mode_o -> rmap_mem_nfee_comm_1:channel_hk_err_invalid_ccd_mode_i
	wire   [15:0] comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_frame_counter_signal;                     // COMM_Pedreiro_v1_01_1:channel_hk_frame_counter_o -> rmap_mem_nfee_comm_1:channel_hk_frame_counter_i
	wire    [1:0] comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_timecode_control_signal;                  // COMM_Pedreiro_v1_01_1:channel_hk_timecode_control_o -> rmap_mem_nfee_comm_1:channel_hk_timecode_control_i
	wire    [1:0] comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_frame_number_signal;                      // COMM_Pedreiro_v1_01_1:channel_hk_frame_number_o -> rmap_mem_nfee_comm_1:channel_hk_frame_number_i
	wire          comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_e_side_buffer_full_signal;            // COMM_Pedreiro_v1_01_2:channel_hk_err_e_side_buffer_full_o -> rmap_mem_nfee_comm_2:channel_hk_err_e_side_buffer_full_i
	wire          comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_escape_err_signal;               // COMM_Pedreiro_v1_01_2:channel_hk_spw_link_escape_err_o -> rmap_mem_nfee_comm_2:channel_hk_spw_link_escape_err_i
	wire          comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_rmap_target_indicate_signal;              // COMM_Pedreiro_v1_01_2:channel_hk_rmap_target_indicate_o -> rmap_mem_nfee_comm_2:channel_hk_rmap_target_indicate_i
	wire          comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal;             // COMM_Pedreiro_v1_01_2:channel_hk_err_win_wrong_y_coord_o -> rmap_mem_nfee_comm_2:channel_hk_err_win_wrong_y_coord_i
	wire          comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_running_signal;                  // COMM_Pedreiro_v1_01_2:channel_hk_spw_link_running_o -> rmap_mem_nfee_comm_2:channel_hk_spw_link_running_i
	wire          comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_credit_err_signal;               // COMM_Pedreiro_v1_01_2:channel_hk_spw_link_credit_err_o -> rmap_mem_nfee_comm_2:channel_hk_spw_link_credit_err_i
	wire          comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal;             // COMM_Pedreiro_v1_01_2:channel_hk_err_win_wrong_x_coord_o -> rmap_mem_nfee_comm_2:channel_hk_err_win_wrong_x_coord_i
	wire    [7:0] comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_rmap_target_status_signal;                // COMM_Pedreiro_v1_01_2:channel_hk_rmap_target_status_o -> rmap_mem_nfee_comm_2:channel_hk_rmap_target_status_i
	wire          comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_f_side_buffer_full_signal;            // COMM_Pedreiro_v1_01_2:channel_hk_err_f_side_buffer_full_o -> rmap_mem_nfee_comm_2:channel_hk_err_f_side_buffer_full_i
	wire    [5:0] comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_timecode_time_signal;                     // COMM_Pedreiro_v1_01_2:channel_hk_timecode_time_o -> rmap_mem_nfee_comm_2:channel_hk_timecode_time_i
	wire          comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_parity_err_signal;               // COMM_Pedreiro_v1_01_2:channel_hk_spw_link_parity_err_o -> rmap_mem_nfee_comm_2:channel_hk_spw_link_parity_err_i
	wire          comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_disconnect_signal;               // COMM_Pedreiro_v1_01_2:channel_hk_spw_link_disconnect_o -> rmap_mem_nfee_comm_2:channel_hk_spw_link_disconnect_i
	wire          comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal;              // COMM_Pedreiro_v1_01_2:channel_hk_err_invalid_ccd_mode_o -> rmap_mem_nfee_comm_2:channel_hk_err_invalid_ccd_mode_i
	wire   [15:0] comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_frame_counter_signal;                     // COMM_Pedreiro_v1_01_2:channel_hk_frame_counter_o -> rmap_mem_nfee_comm_2:channel_hk_frame_counter_i
	wire    [1:0] comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_timecode_control_signal;                  // COMM_Pedreiro_v1_01_2:channel_hk_timecode_control_o -> rmap_mem_nfee_comm_2:channel_hk_timecode_control_i
	wire    [1:0] comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_frame_number_signal;                      // COMM_Pedreiro_v1_01_2:channel_hk_frame_number_o -> rmap_mem_nfee_comm_2:channel_hk_frame_number_i
	wire          comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_e_side_buffer_full_signal;            // COMM_Pedreiro_v1_01_3:channel_hk_err_e_side_buffer_full_o -> rmap_mem_nfee_comm_3:channel_hk_err_e_side_buffer_full_i
	wire          comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_escape_err_signal;               // COMM_Pedreiro_v1_01_3:channel_hk_spw_link_escape_err_o -> rmap_mem_nfee_comm_3:channel_hk_spw_link_escape_err_i
	wire          comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_rmap_target_indicate_signal;              // COMM_Pedreiro_v1_01_3:channel_hk_rmap_target_indicate_o -> rmap_mem_nfee_comm_3:channel_hk_rmap_target_indicate_i
	wire          comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal;             // COMM_Pedreiro_v1_01_3:channel_hk_err_win_wrong_y_coord_o -> rmap_mem_nfee_comm_3:channel_hk_err_win_wrong_y_coord_i
	wire          comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_running_signal;                  // COMM_Pedreiro_v1_01_3:channel_hk_spw_link_running_o -> rmap_mem_nfee_comm_3:channel_hk_spw_link_running_i
	wire          comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_credit_err_signal;               // COMM_Pedreiro_v1_01_3:channel_hk_spw_link_credit_err_o -> rmap_mem_nfee_comm_3:channel_hk_spw_link_credit_err_i
	wire          comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal;             // COMM_Pedreiro_v1_01_3:channel_hk_err_win_wrong_x_coord_o -> rmap_mem_nfee_comm_3:channel_hk_err_win_wrong_x_coord_i
	wire    [7:0] comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_rmap_target_status_signal;                // COMM_Pedreiro_v1_01_3:channel_hk_rmap_target_status_o -> rmap_mem_nfee_comm_3:channel_hk_rmap_target_status_i
	wire          comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_f_side_buffer_full_signal;            // COMM_Pedreiro_v1_01_3:channel_hk_err_f_side_buffer_full_o -> rmap_mem_nfee_comm_3:channel_hk_err_f_side_buffer_full_i
	wire    [5:0] comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_timecode_time_signal;                     // COMM_Pedreiro_v1_01_3:channel_hk_timecode_time_o -> rmap_mem_nfee_comm_3:channel_hk_timecode_time_i
	wire          comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_parity_err_signal;               // COMM_Pedreiro_v1_01_3:channel_hk_spw_link_parity_err_o -> rmap_mem_nfee_comm_3:channel_hk_spw_link_parity_err_i
	wire          comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_disconnect_signal;               // COMM_Pedreiro_v1_01_3:channel_hk_spw_link_disconnect_o -> rmap_mem_nfee_comm_3:channel_hk_spw_link_disconnect_i
	wire          comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal;              // COMM_Pedreiro_v1_01_3:channel_hk_err_invalid_ccd_mode_o -> rmap_mem_nfee_comm_3:channel_hk_err_invalid_ccd_mode_i
	wire   [15:0] comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_frame_counter_signal;                     // COMM_Pedreiro_v1_01_3:channel_hk_frame_counter_o -> rmap_mem_nfee_comm_3:channel_hk_frame_counter_i
	wire    [1:0] comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_timecode_control_signal;                  // COMM_Pedreiro_v1_01_3:channel_hk_timecode_control_o -> rmap_mem_nfee_comm_3:channel_hk_timecode_control_i
	wire    [1:0] comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_frame_number_signal;                      // COMM_Pedreiro_v1_01_3:channel_hk_frame_number_o -> rmap_mem_nfee_comm_3:channel_hk_frame_number_i
	wire          comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_e_side_buffer_full_signal;            // COMM_Pedreiro_v1_01_4:channel_hk_err_e_side_buffer_full_o -> rmap_mem_nfee_comm_4:channel_hk_err_e_side_buffer_full_i
	wire          comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_escape_err_signal;               // COMM_Pedreiro_v1_01_4:channel_hk_spw_link_escape_err_o -> rmap_mem_nfee_comm_4:channel_hk_spw_link_escape_err_i
	wire          comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_rmap_target_indicate_signal;              // COMM_Pedreiro_v1_01_4:channel_hk_rmap_target_indicate_o -> rmap_mem_nfee_comm_4:channel_hk_rmap_target_indicate_i
	wire          comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal;             // COMM_Pedreiro_v1_01_4:channel_hk_err_win_wrong_y_coord_o -> rmap_mem_nfee_comm_4:channel_hk_err_win_wrong_y_coord_i
	wire          comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_running_signal;                  // COMM_Pedreiro_v1_01_4:channel_hk_spw_link_running_o -> rmap_mem_nfee_comm_4:channel_hk_spw_link_running_i
	wire          comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_credit_err_signal;               // COMM_Pedreiro_v1_01_4:channel_hk_spw_link_credit_err_o -> rmap_mem_nfee_comm_4:channel_hk_spw_link_credit_err_i
	wire          comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal;             // COMM_Pedreiro_v1_01_4:channel_hk_err_win_wrong_x_coord_o -> rmap_mem_nfee_comm_4:channel_hk_err_win_wrong_x_coord_i
	wire    [7:0] comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_rmap_target_status_signal;                // COMM_Pedreiro_v1_01_4:channel_hk_rmap_target_status_o -> rmap_mem_nfee_comm_4:channel_hk_rmap_target_status_i
	wire          comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_f_side_buffer_full_signal;            // COMM_Pedreiro_v1_01_4:channel_hk_err_f_side_buffer_full_o -> rmap_mem_nfee_comm_4:channel_hk_err_f_side_buffer_full_i
	wire    [5:0] comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_timecode_time_signal;                     // COMM_Pedreiro_v1_01_4:channel_hk_timecode_time_o -> rmap_mem_nfee_comm_4:channel_hk_timecode_time_i
	wire          comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_parity_err_signal;               // COMM_Pedreiro_v1_01_4:channel_hk_spw_link_parity_err_o -> rmap_mem_nfee_comm_4:channel_hk_spw_link_parity_err_i
	wire          comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_disconnect_signal;               // COMM_Pedreiro_v1_01_4:channel_hk_spw_link_disconnect_o -> rmap_mem_nfee_comm_4:channel_hk_spw_link_disconnect_i
	wire          comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal;              // COMM_Pedreiro_v1_01_4:channel_hk_err_invalid_ccd_mode_o -> rmap_mem_nfee_comm_4:channel_hk_err_invalid_ccd_mode_i
	wire   [15:0] comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_frame_counter_signal;                     // COMM_Pedreiro_v1_01_4:channel_hk_frame_counter_o -> rmap_mem_nfee_comm_4:channel_hk_frame_counter_i
	wire    [1:0] comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_timecode_control_signal;                  // COMM_Pedreiro_v1_01_4:channel_hk_timecode_control_o -> rmap_mem_nfee_comm_4:channel_hk_timecode_control_i
	wire    [1:0] comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_frame_number_signal;                      // COMM_Pedreiro_v1_01_4:channel_hk_frame_number_o -> rmap_mem_nfee_comm_4:channel_hk_frame_number_i
	wire          comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_e_side_buffer_full_signal;            // COMM_Pedreiro_v1_01_6:channel_hk_err_e_side_buffer_full_o -> rmap_mem_nfee_comm_6:channel_hk_err_e_side_buffer_full_i
	wire          comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_escape_err_signal;               // COMM_Pedreiro_v1_01_6:channel_hk_spw_link_escape_err_o -> rmap_mem_nfee_comm_6:channel_hk_spw_link_escape_err_i
	wire          comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_rmap_target_indicate_signal;              // COMM_Pedreiro_v1_01_6:channel_hk_rmap_target_indicate_o -> rmap_mem_nfee_comm_6:channel_hk_rmap_target_indicate_i
	wire          comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal;             // COMM_Pedreiro_v1_01_6:channel_hk_err_win_wrong_y_coord_o -> rmap_mem_nfee_comm_6:channel_hk_err_win_wrong_y_coord_i
	wire          comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_running_signal;                  // COMM_Pedreiro_v1_01_6:channel_hk_spw_link_running_o -> rmap_mem_nfee_comm_6:channel_hk_spw_link_running_i
	wire          comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_credit_err_signal;               // COMM_Pedreiro_v1_01_6:channel_hk_spw_link_credit_err_o -> rmap_mem_nfee_comm_6:channel_hk_spw_link_credit_err_i
	wire          comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal;             // COMM_Pedreiro_v1_01_6:channel_hk_err_win_wrong_x_coord_o -> rmap_mem_nfee_comm_6:channel_hk_err_win_wrong_x_coord_i
	wire    [7:0] comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_rmap_target_status_signal;                // COMM_Pedreiro_v1_01_6:channel_hk_rmap_target_status_o -> rmap_mem_nfee_comm_6:channel_hk_rmap_target_status_i
	wire          comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_f_side_buffer_full_signal;            // COMM_Pedreiro_v1_01_6:channel_hk_err_f_side_buffer_full_o -> rmap_mem_nfee_comm_6:channel_hk_err_f_side_buffer_full_i
	wire    [5:0] comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_timecode_time_signal;                     // COMM_Pedreiro_v1_01_6:channel_hk_timecode_time_o -> rmap_mem_nfee_comm_6:channel_hk_timecode_time_i
	wire          comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_parity_err_signal;               // COMM_Pedreiro_v1_01_6:channel_hk_spw_link_parity_err_o -> rmap_mem_nfee_comm_6:channel_hk_spw_link_parity_err_i
	wire          comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_disconnect_signal;               // COMM_Pedreiro_v1_01_6:channel_hk_spw_link_disconnect_o -> rmap_mem_nfee_comm_6:channel_hk_spw_link_disconnect_i
	wire          comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal;              // COMM_Pedreiro_v1_01_6:channel_hk_err_invalid_ccd_mode_o -> rmap_mem_nfee_comm_6:channel_hk_err_invalid_ccd_mode_i
	wire   [15:0] comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_frame_counter_signal;                     // COMM_Pedreiro_v1_01_6:channel_hk_frame_counter_o -> rmap_mem_nfee_comm_6:channel_hk_frame_counter_i
	wire    [1:0] comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_timecode_control_signal;                  // COMM_Pedreiro_v1_01_6:channel_hk_timecode_control_o -> rmap_mem_nfee_comm_6:channel_hk_timecode_control_i
	wire    [1:0] comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_frame_number_signal;                      // COMM_Pedreiro_v1_01_6:channel_hk_frame_number_o -> rmap_mem_nfee_comm_6:channel_hk_frame_number_i
	wire          comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_e_side_buffer_full_signal;            // COMM_Pedreiro_v1_01_5:channel_hk_err_e_side_buffer_full_o -> rmap_mem_nfee_comm_5:channel_hk_err_e_side_buffer_full_i
	wire          comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_escape_err_signal;               // COMM_Pedreiro_v1_01_5:channel_hk_spw_link_escape_err_o -> rmap_mem_nfee_comm_5:channel_hk_spw_link_escape_err_i
	wire          comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_rmap_target_indicate_signal;              // COMM_Pedreiro_v1_01_5:channel_hk_rmap_target_indicate_o -> rmap_mem_nfee_comm_5:channel_hk_rmap_target_indicate_i
	wire          comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal;             // COMM_Pedreiro_v1_01_5:channel_hk_err_win_wrong_y_coord_o -> rmap_mem_nfee_comm_5:channel_hk_err_win_wrong_y_coord_i
	wire          comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_running_signal;                  // COMM_Pedreiro_v1_01_5:channel_hk_spw_link_running_o -> rmap_mem_nfee_comm_5:channel_hk_spw_link_running_i
	wire          comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_credit_err_signal;               // COMM_Pedreiro_v1_01_5:channel_hk_spw_link_credit_err_o -> rmap_mem_nfee_comm_5:channel_hk_spw_link_credit_err_i
	wire          comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal;             // COMM_Pedreiro_v1_01_5:channel_hk_err_win_wrong_x_coord_o -> rmap_mem_nfee_comm_5:channel_hk_err_win_wrong_x_coord_i
	wire    [7:0] comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_rmap_target_status_signal;                // COMM_Pedreiro_v1_01_5:channel_hk_rmap_target_status_o -> rmap_mem_nfee_comm_5:channel_hk_rmap_target_status_i
	wire          comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_f_side_buffer_full_signal;            // COMM_Pedreiro_v1_01_5:channel_hk_err_f_side_buffer_full_o -> rmap_mem_nfee_comm_5:channel_hk_err_f_side_buffer_full_i
	wire    [5:0] comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_timecode_time_signal;                     // COMM_Pedreiro_v1_01_5:channel_hk_timecode_time_o -> rmap_mem_nfee_comm_5:channel_hk_timecode_time_i
	wire          comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_parity_err_signal;               // COMM_Pedreiro_v1_01_5:channel_hk_spw_link_parity_err_o -> rmap_mem_nfee_comm_5:channel_hk_spw_link_parity_err_i
	wire          comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_disconnect_signal;               // COMM_Pedreiro_v1_01_5:channel_hk_spw_link_disconnect_o -> rmap_mem_nfee_comm_5:channel_hk_spw_link_disconnect_i
	wire          comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal;              // COMM_Pedreiro_v1_01_5:channel_hk_err_invalid_ccd_mode_o -> rmap_mem_nfee_comm_5:channel_hk_err_invalid_ccd_mode_i
	wire   [15:0] comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_frame_counter_signal;                     // COMM_Pedreiro_v1_01_5:channel_hk_frame_counter_o -> rmap_mem_nfee_comm_5:channel_hk_frame_counter_i
	wire    [1:0] comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_timecode_control_signal;                  // COMM_Pedreiro_v1_01_5:channel_hk_timecode_control_o -> rmap_mem_nfee_comm_5:channel_hk_timecode_control_i
	wire    [1:0] comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_frame_number_signal;                      // COMM_Pedreiro_v1_01_5:channel_hk_frame_number_o -> rmap_mem_nfee_comm_5:channel_hk_frame_number_i
	wire          comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_echo_id_en_signal;                     // COMM_Pedreiro_v1_01_1:fee_rmap_echo_id_en_o -> RMAP_Echoing_0:fee_0_rmap_echo_id_en_i
	wire          comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal;      // COMM_Pedreiro_v1_01_1:fee_rmap_incoming_fifo_wrdata_flag_o -> RMAP_Echoing_0:fee_0_rmap_incoming_fifo_wrdata_flag_i
	wire    [7:0] comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal;      // COMM_Pedreiro_v1_01_1:fee_rmap_incoming_fifo_wrdata_data_o -> RMAP_Echoing_0:fee_0_rmap_incoming_fifo_wrdata_data_i
	wire          comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal;            // COMM_Pedreiro_v1_01_1:fee_rmap_incoming_fifo_wrreq_o -> RMAP_Echoing_0:fee_0_rmap_incoming_fifo_wrreq_i
	wire    [7:0] comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal;      // COMM_Pedreiro_v1_01_1:fee_rmap_outgoing_fifo_wrdata_data_o -> RMAP_Echoing_0:fee_0_rmap_outgoing_fifo_wrdata_data_i
	wire          comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal;      // COMM_Pedreiro_v1_01_1:fee_rmap_outgoing_fifo_wrdata_flag_o -> RMAP_Echoing_0:fee_0_rmap_outgoing_fifo_wrdata_flag_i
	wire          comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal;            // COMM_Pedreiro_v1_01_1:fee_rmap_outgoing_fifo_wrreq_o -> RMAP_Echoing_0:fee_0_rmap_outgoing_fifo_wrreq_i
	wire          comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_echo_en_signal;                        // COMM_Pedreiro_v1_01_1:fee_rmap_echo_en_o -> RMAP_Echoing_0:fee_0_rmap_echo_en_i
	wire          comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_echo_id_en_signal;                     // COMM_Pedreiro_v1_01_2:fee_rmap_echo_id_en_o -> RMAP_Echoing_0:fee_1_rmap_echo_id_en_i
	wire          comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal;      // COMM_Pedreiro_v1_01_2:fee_rmap_incoming_fifo_wrdata_flag_o -> RMAP_Echoing_0:fee_1_rmap_incoming_fifo_wrdata_flag_i
	wire    [7:0] comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal;      // COMM_Pedreiro_v1_01_2:fee_rmap_incoming_fifo_wrdata_data_o -> RMAP_Echoing_0:fee_1_rmap_incoming_fifo_wrdata_data_i
	wire          comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal;            // COMM_Pedreiro_v1_01_2:fee_rmap_incoming_fifo_wrreq_o -> RMAP_Echoing_0:fee_1_rmap_incoming_fifo_wrreq_i
	wire    [7:0] comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal;      // COMM_Pedreiro_v1_01_2:fee_rmap_outgoing_fifo_wrdata_data_o -> RMAP_Echoing_0:fee_1_rmap_outgoing_fifo_wrdata_data_i
	wire          comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal;      // COMM_Pedreiro_v1_01_2:fee_rmap_outgoing_fifo_wrdata_flag_o -> RMAP_Echoing_0:fee_1_rmap_outgoing_fifo_wrdata_flag_i
	wire          comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal;            // COMM_Pedreiro_v1_01_2:fee_rmap_outgoing_fifo_wrreq_o -> RMAP_Echoing_0:fee_1_rmap_outgoing_fifo_wrreq_i
	wire          comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_echo_en_signal;                        // COMM_Pedreiro_v1_01_2:fee_rmap_echo_en_o -> RMAP_Echoing_0:fee_1_rmap_echo_en_i
	wire          comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_echo_id_en_signal;                     // COMM_Pedreiro_v1_01_4:fee_rmap_echo_id_en_o -> RMAP_Echoing_0:fee_3_rmap_echo_id_en_i
	wire          comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal;      // COMM_Pedreiro_v1_01_4:fee_rmap_incoming_fifo_wrdata_flag_o -> RMAP_Echoing_0:fee_3_rmap_incoming_fifo_wrdata_flag_i
	wire    [7:0] comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal;      // COMM_Pedreiro_v1_01_4:fee_rmap_incoming_fifo_wrdata_data_o -> RMAP_Echoing_0:fee_3_rmap_incoming_fifo_wrdata_data_i
	wire          comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal;            // COMM_Pedreiro_v1_01_4:fee_rmap_incoming_fifo_wrreq_o -> RMAP_Echoing_0:fee_3_rmap_incoming_fifo_wrreq_i
	wire    [7:0] comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal;      // COMM_Pedreiro_v1_01_4:fee_rmap_outgoing_fifo_wrdata_data_o -> RMAP_Echoing_0:fee_3_rmap_outgoing_fifo_wrdata_data_i
	wire          comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal;      // COMM_Pedreiro_v1_01_4:fee_rmap_outgoing_fifo_wrdata_flag_o -> RMAP_Echoing_0:fee_3_rmap_outgoing_fifo_wrdata_flag_i
	wire          comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal;            // COMM_Pedreiro_v1_01_4:fee_rmap_outgoing_fifo_wrreq_o -> RMAP_Echoing_0:fee_3_rmap_outgoing_fifo_wrreq_i
	wire          comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_echo_en_signal;                        // COMM_Pedreiro_v1_01_4:fee_rmap_echo_en_o -> RMAP_Echoing_0:fee_3_rmap_echo_en_i
	wire          comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_echo_id_en_signal;                     // COMM_Pedreiro_v1_01_5:fee_rmap_echo_id_en_o -> RMAP_Echoing_0:fee_4_rmap_echo_id_en_i
	wire          comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal;      // COMM_Pedreiro_v1_01_5:fee_rmap_incoming_fifo_wrdata_flag_o -> RMAP_Echoing_0:fee_4_rmap_incoming_fifo_wrdata_flag_i
	wire    [7:0] comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal;      // COMM_Pedreiro_v1_01_5:fee_rmap_incoming_fifo_wrdata_data_o -> RMAP_Echoing_0:fee_4_rmap_incoming_fifo_wrdata_data_i
	wire          comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal;            // COMM_Pedreiro_v1_01_5:fee_rmap_incoming_fifo_wrreq_o -> RMAP_Echoing_0:fee_4_rmap_incoming_fifo_wrreq_i
	wire    [7:0] comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal;      // COMM_Pedreiro_v1_01_5:fee_rmap_outgoing_fifo_wrdata_data_o -> RMAP_Echoing_0:fee_4_rmap_outgoing_fifo_wrdata_data_i
	wire          comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal;      // COMM_Pedreiro_v1_01_5:fee_rmap_outgoing_fifo_wrdata_flag_o -> RMAP_Echoing_0:fee_4_rmap_outgoing_fifo_wrdata_flag_i
	wire          comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal;            // COMM_Pedreiro_v1_01_5:fee_rmap_outgoing_fifo_wrreq_o -> RMAP_Echoing_0:fee_4_rmap_outgoing_fifo_wrreq_i
	wire          comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_echo_en_signal;                        // COMM_Pedreiro_v1_01_5:fee_rmap_echo_en_o -> RMAP_Echoing_0:fee_4_rmap_echo_en_i
	wire          comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_echo_id_en_signal;                     // COMM_Pedreiro_v1_01_6:fee_rmap_echo_id_en_o -> RMAP_Echoing_0:fee_5_rmap_echo_id_en_i
	wire          comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal;      // COMM_Pedreiro_v1_01_6:fee_rmap_incoming_fifo_wrdata_flag_o -> RMAP_Echoing_0:fee_5_rmap_incoming_fifo_wrdata_flag_i
	wire    [7:0] comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal;      // COMM_Pedreiro_v1_01_6:fee_rmap_incoming_fifo_wrdata_data_o -> RMAP_Echoing_0:fee_5_rmap_incoming_fifo_wrdata_data_i
	wire          comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal;            // COMM_Pedreiro_v1_01_6:fee_rmap_incoming_fifo_wrreq_o -> RMAP_Echoing_0:fee_5_rmap_incoming_fifo_wrreq_i
	wire    [7:0] comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal;      // COMM_Pedreiro_v1_01_6:fee_rmap_outgoing_fifo_wrdata_data_o -> RMAP_Echoing_0:fee_5_rmap_outgoing_fifo_wrdata_data_i
	wire          comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal;      // COMM_Pedreiro_v1_01_6:fee_rmap_outgoing_fifo_wrdata_flag_o -> RMAP_Echoing_0:fee_5_rmap_outgoing_fifo_wrdata_flag_i
	wire          comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal;            // COMM_Pedreiro_v1_01_6:fee_rmap_outgoing_fifo_wrreq_o -> RMAP_Echoing_0:fee_5_rmap_outgoing_fifo_wrreq_i
	wire          comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_echo_en_signal;                        // COMM_Pedreiro_v1_01_6:fee_rmap_echo_en_o -> RMAP_Echoing_0:fee_5_rmap_echo_en_i
	wire          comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_echo_id_en_signal;                     // COMM_Pedreiro_v1_01_3:fee_rmap_echo_id_en_o -> RMAP_Echoing_0:fee_2_rmap_echo_id_en_i
	wire          comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal;      // COMM_Pedreiro_v1_01_3:fee_rmap_incoming_fifo_wrdata_flag_o -> RMAP_Echoing_0:fee_2_rmap_incoming_fifo_wrdata_flag_i
	wire    [7:0] comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal;      // COMM_Pedreiro_v1_01_3:fee_rmap_incoming_fifo_wrdata_data_o -> RMAP_Echoing_0:fee_2_rmap_incoming_fifo_wrdata_data_i
	wire          comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal;            // COMM_Pedreiro_v1_01_3:fee_rmap_incoming_fifo_wrreq_o -> RMAP_Echoing_0:fee_2_rmap_incoming_fifo_wrreq_i
	wire    [7:0] comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal;      // COMM_Pedreiro_v1_01_3:fee_rmap_outgoing_fifo_wrdata_data_o -> RMAP_Echoing_0:fee_2_rmap_outgoing_fifo_wrdata_data_i
	wire          comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal;      // COMM_Pedreiro_v1_01_3:fee_rmap_outgoing_fifo_wrdata_flag_o -> RMAP_Echoing_0:fee_2_rmap_outgoing_fifo_wrdata_flag_i
	wire          comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal;            // COMM_Pedreiro_v1_01_3:fee_rmap_outgoing_fifo_wrreq_o -> RMAP_Echoing_0:fee_2_rmap_outgoing_fifo_wrreq_i
	wire          comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_echo_en_signal;                        // COMM_Pedreiro_v1_01_3:fee_rmap_echo_en_o -> RMAP_Echoing_0:fee_2_rmap_echo_en_i
	wire          comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_write_signal;                      // COMM_Pedreiro_v1_01_3:fee_codec_rmap_write_o -> rmap_mem_nfee_comm_3:fee_0_rmap_write_i
	wire    [7:0] rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_readdata_signal;                         // rmap_mem_nfee_comm_3:fee_0_rmap_readdata_o -> COMM_Pedreiro_v1_01_3:fee_codec_rmap_readdata_i
	wire   [31:0] comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_rd_address_signal;                 // COMM_Pedreiro_v1_01_3:fee_codec_rmap_rd_address_o -> rmap_mem_nfee_comm_3:fee_0_rmap_rd_address_i
	wire   [31:0] comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_wr_address_signal;                 // COMM_Pedreiro_v1_01_3:fee_codec_rmap_wr_address_o -> rmap_mem_nfee_comm_3:fee_0_rmap_wr_address_i
	wire          comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_read_signal;                       // COMM_Pedreiro_v1_01_3:fee_codec_rmap_read_o -> rmap_mem_nfee_comm_3:fee_0_rmap_read_i
	wire          rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal;                   // rmap_mem_nfee_comm_3:fee_0_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_3:fee_codec_rmap_wr_waitrequest_i
	wire          rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal;                   // rmap_mem_nfee_comm_3:fee_0_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_3:fee_codec_rmap_rd_waitrequest_i
	wire    [7:0] comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_writedata_signal;                  // COMM_Pedreiro_v1_01_3:fee_codec_rmap_writedata_o -> rmap_mem_nfee_comm_3:fee_0_rmap_writedata_i
	wire          comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_write_signal;                      // COMM_Pedreiro_v1_01_1:fee_codec_rmap_write_o -> rmap_mem_nfee_comm_1:fee_0_rmap_write_i
	wire   [31:0] comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_rd_address_signal;                 // COMM_Pedreiro_v1_01_1:fee_codec_rmap_rd_address_o -> rmap_mem_nfee_comm_1:fee_0_rmap_rd_address_i
	wire    [7:0] rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_readdata_signal;                         // rmap_mem_nfee_comm_1:fee_0_rmap_readdata_o -> COMM_Pedreiro_v1_01_1:fee_codec_rmap_readdata_i
	wire   [31:0] comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_wr_address_signal;                 // COMM_Pedreiro_v1_01_1:fee_codec_rmap_wr_address_o -> rmap_mem_nfee_comm_1:fee_0_rmap_wr_address_i
	wire          comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_read_signal;                       // COMM_Pedreiro_v1_01_1:fee_codec_rmap_read_o -> rmap_mem_nfee_comm_1:fee_0_rmap_read_i
	wire          rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal;                   // rmap_mem_nfee_comm_1:fee_0_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_1:fee_codec_rmap_wr_waitrequest_i
	wire    [7:0] comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_writedata_signal;                  // COMM_Pedreiro_v1_01_1:fee_codec_rmap_writedata_o -> rmap_mem_nfee_comm_1:fee_0_rmap_writedata_i
	wire          rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal;                   // rmap_mem_nfee_comm_1:fee_0_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_1:fee_codec_rmap_rd_waitrequest_i
	wire          comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_write_signal;                      // COMM_Pedreiro_v1_01_2:fee_codec_rmap_write_o -> rmap_mem_nfee_comm_2:fee_0_rmap_write_i
	wire   [31:0] comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_rd_address_signal;                 // COMM_Pedreiro_v1_01_2:fee_codec_rmap_rd_address_o -> rmap_mem_nfee_comm_2:fee_0_rmap_rd_address_i
	wire    [7:0] rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_readdata_signal;                         // rmap_mem_nfee_comm_2:fee_0_rmap_readdata_o -> COMM_Pedreiro_v1_01_2:fee_codec_rmap_readdata_i
	wire   [31:0] comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_wr_address_signal;                 // COMM_Pedreiro_v1_01_2:fee_codec_rmap_wr_address_o -> rmap_mem_nfee_comm_2:fee_0_rmap_wr_address_i
	wire          comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_read_signal;                       // COMM_Pedreiro_v1_01_2:fee_codec_rmap_read_o -> rmap_mem_nfee_comm_2:fee_0_rmap_read_i
	wire          rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal;                   // rmap_mem_nfee_comm_2:fee_0_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_2:fee_codec_rmap_wr_waitrequest_i
	wire    [7:0] comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_writedata_signal;                  // COMM_Pedreiro_v1_01_2:fee_codec_rmap_writedata_o -> rmap_mem_nfee_comm_2:fee_0_rmap_writedata_i
	wire          rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal;                   // rmap_mem_nfee_comm_2:fee_0_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_2:fee_codec_rmap_rd_waitrequest_i
	wire          comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_write_signal;                      // COMM_Pedreiro_v1_01_4:fee_codec_rmap_write_o -> rmap_mem_nfee_comm_4:fee_0_rmap_write_i
	wire   [31:0] comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_rd_address_signal;                 // COMM_Pedreiro_v1_01_4:fee_codec_rmap_rd_address_o -> rmap_mem_nfee_comm_4:fee_0_rmap_rd_address_i
	wire    [7:0] rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_readdata_signal;                         // rmap_mem_nfee_comm_4:fee_0_rmap_readdata_o -> COMM_Pedreiro_v1_01_4:fee_codec_rmap_readdata_i
	wire   [31:0] comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_wr_address_signal;                 // COMM_Pedreiro_v1_01_4:fee_codec_rmap_wr_address_o -> rmap_mem_nfee_comm_4:fee_0_rmap_wr_address_i
	wire          comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_read_signal;                       // COMM_Pedreiro_v1_01_4:fee_codec_rmap_read_o -> rmap_mem_nfee_comm_4:fee_0_rmap_read_i
	wire          rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal;                   // rmap_mem_nfee_comm_4:fee_0_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_4:fee_codec_rmap_wr_waitrequest_i
	wire    [7:0] comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_writedata_signal;                  // COMM_Pedreiro_v1_01_4:fee_codec_rmap_writedata_o -> rmap_mem_nfee_comm_4:fee_0_rmap_writedata_i
	wire          rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal;                   // rmap_mem_nfee_comm_4:fee_0_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_4:fee_codec_rmap_rd_waitrequest_i
	wire          comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_write_signal;                      // COMM_Pedreiro_v1_01_5:fee_codec_rmap_write_o -> rmap_mem_nfee_comm_5:fee_0_rmap_write_i
	wire   [31:0] comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_rd_address_signal;                 // COMM_Pedreiro_v1_01_5:fee_codec_rmap_rd_address_o -> rmap_mem_nfee_comm_5:fee_0_rmap_rd_address_i
	wire    [7:0] rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_readdata_signal;                         // rmap_mem_nfee_comm_5:fee_0_rmap_readdata_o -> COMM_Pedreiro_v1_01_5:fee_codec_rmap_readdata_i
	wire   [31:0] comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_wr_address_signal;                 // COMM_Pedreiro_v1_01_5:fee_codec_rmap_wr_address_o -> rmap_mem_nfee_comm_5:fee_0_rmap_wr_address_i
	wire          comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_read_signal;                       // COMM_Pedreiro_v1_01_5:fee_codec_rmap_read_o -> rmap_mem_nfee_comm_5:fee_0_rmap_read_i
	wire          rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal;                   // rmap_mem_nfee_comm_5:fee_0_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_5:fee_codec_rmap_wr_waitrequest_i
	wire    [7:0] comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_writedata_signal;                  // COMM_Pedreiro_v1_01_5:fee_codec_rmap_writedata_o -> rmap_mem_nfee_comm_5:fee_0_rmap_writedata_i
	wire          rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal;                   // rmap_mem_nfee_comm_5:fee_0_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_5:fee_codec_rmap_rd_waitrequest_i
	wire          comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_write_signal;                      // COMM_Pedreiro_v1_01_6:fee_codec_rmap_write_o -> rmap_mem_nfee_comm_6:fee_0_rmap_write_i
	wire   [31:0] comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_rd_address_signal;                 // COMM_Pedreiro_v1_01_6:fee_codec_rmap_rd_address_o -> rmap_mem_nfee_comm_6:fee_0_rmap_rd_address_i
	wire    [7:0] rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_readdata_signal;                         // rmap_mem_nfee_comm_6:fee_0_rmap_readdata_o -> COMM_Pedreiro_v1_01_6:fee_codec_rmap_readdata_i
	wire   [31:0] comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_wr_address_signal;                 // COMM_Pedreiro_v1_01_6:fee_codec_rmap_wr_address_o -> rmap_mem_nfee_comm_6:fee_0_rmap_wr_address_i
	wire          comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_read_signal;                       // COMM_Pedreiro_v1_01_6:fee_codec_rmap_read_o -> rmap_mem_nfee_comm_6:fee_0_rmap_read_i
	wire          rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal;                   // rmap_mem_nfee_comm_6:fee_0_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_6:fee_codec_rmap_wr_waitrequest_i
	wire    [7:0] comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_writedata_signal;                  // COMM_Pedreiro_v1_01_6:fee_codec_rmap_writedata_o -> rmap_mem_nfee_comm_6:fee_0_rmap_writedata_i
	wire          rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal;                   // rmap_mem_nfee_comm_6:fee_0_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_6:fee_codec_rmap_rd_waitrequest_i
	wire          comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_write_signal;                         // COMM_Pedreiro_v1_01_1:fee_hk_rmap_write_o -> rmap_mem_nfee_comm_1:fee_1_rmap_write_i
	wire   [31:0] comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_rd_address_signal;                    // COMM_Pedreiro_v1_01_1:fee_hk_rmap_rd_address_o -> rmap_mem_nfee_comm_1:fee_1_rmap_rd_address_i
	wire    [7:0] rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_readdata_signal;                         // rmap_mem_nfee_comm_1:fee_1_rmap_readdata_o -> COMM_Pedreiro_v1_01_1:fee_hk_rmap_readdata_i
	wire   [31:0] comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_wr_address_signal;                    // COMM_Pedreiro_v1_01_1:fee_hk_rmap_wr_address_o -> rmap_mem_nfee_comm_1:fee_1_rmap_wr_address_i
	wire          comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_read_signal;                          // COMM_Pedreiro_v1_01_1:fee_hk_rmap_read_o -> rmap_mem_nfee_comm_1:fee_1_rmap_read_i
	wire          rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal;                   // rmap_mem_nfee_comm_1:fee_1_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_1:fee_hk_rmap_wr_waitrequest_i
	wire    [7:0] comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_writedata_signal;                     // COMM_Pedreiro_v1_01_1:fee_hk_rmap_writedata_o -> rmap_mem_nfee_comm_1:fee_1_rmap_writedata_i
	wire          rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal;                   // rmap_mem_nfee_comm_1:fee_1_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_1:fee_hk_rmap_rd_waitrequest_i
	wire          comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_write_signal;                         // COMM_Pedreiro_v1_01_2:fee_hk_rmap_write_o -> rmap_mem_nfee_comm_2:fee_1_rmap_write_i
	wire   [31:0] comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_rd_address_signal;                    // COMM_Pedreiro_v1_01_2:fee_hk_rmap_rd_address_o -> rmap_mem_nfee_comm_2:fee_1_rmap_rd_address_i
	wire    [7:0] rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_readdata_signal;                         // rmap_mem_nfee_comm_2:fee_1_rmap_readdata_o -> COMM_Pedreiro_v1_01_2:fee_hk_rmap_readdata_i
	wire   [31:0] comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_wr_address_signal;                    // COMM_Pedreiro_v1_01_2:fee_hk_rmap_wr_address_o -> rmap_mem_nfee_comm_2:fee_1_rmap_wr_address_i
	wire          comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_read_signal;                          // COMM_Pedreiro_v1_01_2:fee_hk_rmap_read_o -> rmap_mem_nfee_comm_2:fee_1_rmap_read_i
	wire          rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal;                   // rmap_mem_nfee_comm_2:fee_1_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_2:fee_hk_rmap_wr_waitrequest_i
	wire    [7:0] comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_writedata_signal;                     // COMM_Pedreiro_v1_01_2:fee_hk_rmap_writedata_o -> rmap_mem_nfee_comm_2:fee_1_rmap_writedata_i
	wire          rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal;                   // rmap_mem_nfee_comm_2:fee_1_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_2:fee_hk_rmap_rd_waitrequest_i
	wire          comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_write_signal;                         // COMM_Pedreiro_v1_01_3:fee_hk_rmap_write_o -> rmap_mem_nfee_comm_3:fee_1_rmap_write_i
	wire   [31:0] comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_rd_address_signal;                    // COMM_Pedreiro_v1_01_3:fee_hk_rmap_rd_address_o -> rmap_mem_nfee_comm_3:fee_1_rmap_rd_address_i
	wire    [7:0] rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_readdata_signal;                         // rmap_mem_nfee_comm_3:fee_1_rmap_readdata_o -> COMM_Pedreiro_v1_01_3:fee_hk_rmap_readdata_i
	wire   [31:0] comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_wr_address_signal;                    // COMM_Pedreiro_v1_01_3:fee_hk_rmap_wr_address_o -> rmap_mem_nfee_comm_3:fee_1_rmap_wr_address_i
	wire          comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_read_signal;                          // COMM_Pedreiro_v1_01_3:fee_hk_rmap_read_o -> rmap_mem_nfee_comm_3:fee_1_rmap_read_i
	wire          rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal;                   // rmap_mem_nfee_comm_3:fee_1_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_3:fee_hk_rmap_wr_waitrequest_i
	wire    [7:0] comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_writedata_signal;                     // COMM_Pedreiro_v1_01_3:fee_hk_rmap_writedata_o -> rmap_mem_nfee_comm_3:fee_1_rmap_writedata_i
	wire          rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal;                   // rmap_mem_nfee_comm_3:fee_1_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_3:fee_hk_rmap_rd_waitrequest_i
	wire          comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_write_signal;                         // COMM_Pedreiro_v1_01_4:fee_hk_rmap_write_o -> rmap_mem_nfee_comm_4:fee_1_rmap_write_i
	wire   [31:0] comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_rd_address_signal;                    // COMM_Pedreiro_v1_01_4:fee_hk_rmap_rd_address_o -> rmap_mem_nfee_comm_4:fee_1_rmap_rd_address_i
	wire    [7:0] rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_readdata_signal;                         // rmap_mem_nfee_comm_4:fee_1_rmap_readdata_o -> COMM_Pedreiro_v1_01_4:fee_hk_rmap_readdata_i
	wire   [31:0] comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_wr_address_signal;                    // COMM_Pedreiro_v1_01_4:fee_hk_rmap_wr_address_o -> rmap_mem_nfee_comm_4:fee_1_rmap_wr_address_i
	wire          comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_read_signal;                          // COMM_Pedreiro_v1_01_4:fee_hk_rmap_read_o -> rmap_mem_nfee_comm_4:fee_1_rmap_read_i
	wire          rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal;                   // rmap_mem_nfee_comm_4:fee_1_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_4:fee_hk_rmap_wr_waitrequest_i
	wire    [7:0] comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_writedata_signal;                     // COMM_Pedreiro_v1_01_4:fee_hk_rmap_writedata_o -> rmap_mem_nfee_comm_4:fee_1_rmap_writedata_i
	wire          rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal;                   // rmap_mem_nfee_comm_4:fee_1_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_4:fee_hk_rmap_rd_waitrequest_i
	wire          comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_write_signal;                         // COMM_Pedreiro_v1_01_5:fee_hk_rmap_write_o -> rmap_mem_nfee_comm_5:fee_1_rmap_write_i
	wire   [31:0] comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_rd_address_signal;                    // COMM_Pedreiro_v1_01_5:fee_hk_rmap_rd_address_o -> rmap_mem_nfee_comm_5:fee_1_rmap_rd_address_i
	wire    [7:0] rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_readdata_signal;                         // rmap_mem_nfee_comm_5:fee_1_rmap_readdata_o -> COMM_Pedreiro_v1_01_5:fee_hk_rmap_readdata_i
	wire   [31:0] comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_wr_address_signal;                    // COMM_Pedreiro_v1_01_5:fee_hk_rmap_wr_address_o -> rmap_mem_nfee_comm_5:fee_1_rmap_wr_address_i
	wire          comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_read_signal;                          // COMM_Pedreiro_v1_01_5:fee_hk_rmap_read_o -> rmap_mem_nfee_comm_5:fee_1_rmap_read_i
	wire          rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal;                   // rmap_mem_nfee_comm_5:fee_1_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_5:fee_hk_rmap_wr_waitrequest_i
	wire    [7:0] comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_writedata_signal;                     // COMM_Pedreiro_v1_01_5:fee_hk_rmap_writedata_o -> rmap_mem_nfee_comm_5:fee_1_rmap_writedata_i
	wire          rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal;                   // rmap_mem_nfee_comm_5:fee_1_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_5:fee_hk_rmap_rd_waitrequest_i
	wire          comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_write_signal;                         // COMM_Pedreiro_v1_01_6:fee_hk_rmap_write_o -> rmap_mem_nfee_comm_6:fee_1_rmap_write_i
	wire   [31:0] comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_rd_address_signal;                    // COMM_Pedreiro_v1_01_6:fee_hk_rmap_rd_address_o -> rmap_mem_nfee_comm_6:fee_1_rmap_rd_address_i
	wire    [7:0] rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_readdata_signal;                         // rmap_mem_nfee_comm_6:fee_1_rmap_readdata_o -> COMM_Pedreiro_v1_01_6:fee_hk_rmap_readdata_i
	wire   [31:0] comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_wr_address_signal;                    // COMM_Pedreiro_v1_01_6:fee_hk_rmap_wr_address_o -> rmap_mem_nfee_comm_6:fee_1_rmap_wr_address_i
	wire          comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_read_signal;                          // COMM_Pedreiro_v1_01_6:fee_hk_rmap_read_o -> rmap_mem_nfee_comm_6:fee_1_rmap_read_i
	wire          rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal;                   // rmap_mem_nfee_comm_6:fee_1_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_6:fee_hk_rmap_wr_waitrequest_i
	wire    [7:0] comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_writedata_signal;                     // COMM_Pedreiro_v1_01_6:fee_hk_rmap_writedata_o -> rmap_mem_nfee_comm_6:fee_1_rmap_writedata_i
	wire          rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal;                   // rmap_mem_nfee_comm_6:fee_1_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_6:fee_hk_rmap_rd_waitrequest_i
	wire   [63:0] comm_pedreiro_v1_01_6_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal;         // COMM_Pedreiro_v1_01_6:channel_win_mem_addr_offset_o -> rmap_mem_nfee_comm_6:channel_win_mem_addr_offset_i
	wire   [63:0] comm_pedreiro_v1_01_1_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal;         // COMM_Pedreiro_v1_01_1:channel_win_mem_addr_offset_o -> rmap_mem_nfee_comm_1:channel_win_mem_addr_offset_i
	wire   [63:0] comm_pedreiro_v1_01_2_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal;         // COMM_Pedreiro_v1_01_2:channel_win_mem_addr_offset_o -> rmap_mem_nfee_comm_2:channel_win_mem_addr_offset_i
	wire   [63:0] comm_pedreiro_v1_01_3_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal;         // COMM_Pedreiro_v1_01_3:channel_win_mem_addr_offset_o -> rmap_mem_nfee_comm_3:channel_win_mem_addr_offset_i
	wire   [63:0] comm_pedreiro_v1_01_4_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal;         // COMM_Pedreiro_v1_01_4:channel_win_mem_addr_offset_o -> rmap_mem_nfee_comm_4:channel_win_mem_addr_offset_i
	wire   [63:0] comm_pedreiro_v1_01_5_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal;         // COMM_Pedreiro_v1_01_5:channel_win_mem_addr_offset_o -> rmap_mem_nfee_comm_5:channel_win_mem_addr_offset_i
	wire          spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal;       // SpaceWire_Channel_A:spw_data_rx_status_rxvalid_o -> COMM_Pedreiro_v1_01_1:spw_data_rx_status_rxvalid_i
	wire    [7:0] comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal;  // COMM_Pedreiro_v1_01_1:spw_data_tx_command_txdata_o -> SpaceWire_Channel_A:spw_data_tx_command_txdata_i
	wire          spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errdisc_signal;           // SpaceWire_Channel_A:spw_link_error_errdisc_o -> COMM_Pedreiro_v1_01_1:spw_link_error_errdisc_i
	wire          spacewire_channel_a_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal;       // SpaceWire_Channel_A:spw_data_tx_status_txhalff_o -> COMM_Pedreiro_v1_01_1:spw_data_tx_status_txhalff_i
	wire          comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal; // COMM_Pedreiro_v1_01_1:spw_data_tx_command_txwrite_o -> SpaceWire_Channel_A:spw_data_tx_command_txwrite_i
	wire          spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal;         // SpaceWire_Channel_A:spw_timecode_rx_tick_out_o -> COMM_Pedreiro_v1_01_1:spw_timecode_rx_tick_out_i
	wire          spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal;       // SpaceWire_Channel_A:spw_data_rx_status_rxhalff_o -> COMM_Pedreiro_v1_01_1:spw_data_rx_status_rxhalff_i
	wire    [5:0] spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal;         // SpaceWire_Channel_A:spw_timecode_rx_time_out_o -> COMM_Pedreiro_v1_01_1:spw_timecode_rx_time_out_i
	wire          spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_connecting_signal;       // SpaceWire_Channel_A:spw_link_status_connecting_o -> COMM_Pedreiro_v1_01_1:spw_link_status_connecting_i
	wire    [7:0] spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal;        // SpaceWire_Channel_A:spw_data_rx_status_rxdata_o -> COMM_Pedreiro_v1_01_1:spw_data_rx_status_rxdata_i
	wire    [1:0] spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal;         // SpaceWire_Channel_A:spw_timecode_rx_ctrl_out_o -> COMM_Pedreiro_v1_01_1:spw_timecode_rx_ctrl_out_i
	wire          comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal;  // COMM_Pedreiro_v1_01_1:spw_data_tx_command_txflag_o -> SpaceWire_Channel_A:spw_data_tx_command_txflag_i
	wire          comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_link_command_linkstart_signal;  // COMM_Pedreiro_v1_01_1:spw_link_command_linkstart_o -> SpaceWire_Channel_A:spw_link_command_linkstart_i
	wire          comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal;  // COMM_Pedreiro_v1_01_1:spw_data_rx_command_rxread_o -> SpaceWire_Channel_A:spw_data_rx_command_rxread_i
	wire          spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_running_signal;          // SpaceWire_Channel_A:spw_link_status_running_o -> COMM_Pedreiro_v1_01_1:spw_link_status_running_i
	wire          spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_started_signal;          // SpaceWire_Channel_A:spw_link_status_started_o -> COMM_Pedreiro_v1_01_1:spw_link_status_started_i
	wire          spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errpar_signal;            // SpaceWire_Channel_A:spw_link_error_errpar_o -> COMM_Pedreiro_v1_01_1:spw_link_error_errpar_i
	wire          comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_link_command_linkdis_signal;    // COMM_Pedreiro_v1_01_1:spw_link_command_linkdis_o -> SpaceWire_Channel_A:spw_link_command_linkdis_i
	wire          spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_erresc_signal;            // SpaceWire_Channel_A:spw_link_error_erresc_o -> COMM_Pedreiro_v1_01_1:spw_link_error_erresc_i
	wire          spacewire_channel_a_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal;         // SpaceWire_Channel_A:spw_data_tx_status_txrdy_o -> COMM_Pedreiro_v1_01_1:spw_data_tx_status_txrdy_i
	wire          comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal;     // COMM_Pedreiro_v1_01_1:spw_timecode_tx_tick_in_o -> SpaceWire_Channel_A:spw_timecode_tx_tick_in_i
	wire    [7:0] comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal;   // COMM_Pedreiro_v1_01_1:spw_link_command_txdivcnt_o -> SpaceWire_Channel_A:spw_link_command_txdivcnt_i
	wire    [5:0] comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal;     // COMM_Pedreiro_v1_01_1:spw_timecode_tx_time_in_o -> SpaceWire_Channel_A:spw_timecode_tx_time_in_i
	wire          spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal;        // SpaceWire_Channel_A:spw_data_rx_status_rxflag_o -> COMM_Pedreiro_v1_01_1:spw_data_rx_status_rxflag_i
	wire    [1:0] comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal;     // COMM_Pedreiro_v1_01_1:spw_timecode_tx_ctrl_in_o -> SpaceWire_Channel_A:spw_timecode_tx_ctrl_in_i
	wire          comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_link_command_autostart_signal;  // COMM_Pedreiro_v1_01_1:spw_link_command_autostart_o -> SpaceWire_Channel_A:spw_link_command_autostart_i
	wire          spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errcred_signal;           // SpaceWire_Channel_A:spw_link_error_errcred_o -> COMM_Pedreiro_v1_01_1:spw_link_error_errcred_i
	wire          spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal;       // SpaceWire_Channel_B:spw_data_rx_status_rxvalid_o -> COMM_Pedreiro_v1_01_2:spw_data_rx_status_rxvalid_i
	wire    [7:0] comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal;  // COMM_Pedreiro_v1_01_2:spw_data_tx_command_txdata_o -> SpaceWire_Channel_B:spw_data_tx_command_txdata_i
	wire          spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errdisc_signal;           // SpaceWire_Channel_B:spw_link_error_errdisc_o -> COMM_Pedreiro_v1_01_2:spw_link_error_errdisc_i
	wire          spacewire_channel_b_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal;       // SpaceWire_Channel_B:spw_data_tx_status_txhalff_o -> COMM_Pedreiro_v1_01_2:spw_data_tx_status_txhalff_i
	wire          comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal; // COMM_Pedreiro_v1_01_2:spw_data_tx_command_txwrite_o -> SpaceWire_Channel_B:spw_data_tx_command_txwrite_i
	wire          spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal;         // SpaceWire_Channel_B:spw_timecode_rx_tick_out_o -> COMM_Pedreiro_v1_01_2:spw_timecode_rx_tick_out_i
	wire          spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal;       // SpaceWire_Channel_B:spw_data_rx_status_rxhalff_o -> COMM_Pedreiro_v1_01_2:spw_data_rx_status_rxhalff_i
	wire    [5:0] spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal;         // SpaceWire_Channel_B:spw_timecode_rx_time_out_o -> COMM_Pedreiro_v1_01_2:spw_timecode_rx_time_out_i
	wire          spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_connecting_signal;       // SpaceWire_Channel_B:spw_link_status_connecting_o -> COMM_Pedreiro_v1_01_2:spw_link_status_connecting_i
	wire    [7:0] spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal;        // SpaceWire_Channel_B:spw_data_rx_status_rxdata_o -> COMM_Pedreiro_v1_01_2:spw_data_rx_status_rxdata_i
	wire    [1:0] spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal;         // SpaceWire_Channel_B:spw_timecode_rx_ctrl_out_o -> COMM_Pedreiro_v1_01_2:spw_timecode_rx_ctrl_out_i
	wire          comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal;  // COMM_Pedreiro_v1_01_2:spw_data_tx_command_txflag_o -> SpaceWire_Channel_B:spw_data_tx_command_txflag_i
	wire          comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_link_command_linkstart_signal;  // COMM_Pedreiro_v1_01_2:spw_link_command_linkstart_o -> SpaceWire_Channel_B:spw_link_command_linkstart_i
	wire          comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal;  // COMM_Pedreiro_v1_01_2:spw_data_rx_command_rxread_o -> SpaceWire_Channel_B:spw_data_rx_command_rxread_i
	wire          spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_running_signal;          // SpaceWire_Channel_B:spw_link_status_running_o -> COMM_Pedreiro_v1_01_2:spw_link_status_running_i
	wire          spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_started_signal;          // SpaceWire_Channel_B:spw_link_status_started_o -> COMM_Pedreiro_v1_01_2:spw_link_status_started_i
	wire          spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errpar_signal;            // SpaceWire_Channel_B:spw_link_error_errpar_o -> COMM_Pedreiro_v1_01_2:spw_link_error_errpar_i
	wire          comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_link_command_linkdis_signal;    // COMM_Pedreiro_v1_01_2:spw_link_command_linkdis_o -> SpaceWire_Channel_B:spw_link_command_linkdis_i
	wire          spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_erresc_signal;            // SpaceWire_Channel_B:spw_link_error_erresc_o -> COMM_Pedreiro_v1_01_2:spw_link_error_erresc_i
	wire          spacewire_channel_b_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal;         // SpaceWire_Channel_B:spw_data_tx_status_txrdy_o -> COMM_Pedreiro_v1_01_2:spw_data_tx_status_txrdy_i
	wire          comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal;     // COMM_Pedreiro_v1_01_2:spw_timecode_tx_tick_in_o -> SpaceWire_Channel_B:spw_timecode_tx_tick_in_i
	wire    [7:0] comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal;   // COMM_Pedreiro_v1_01_2:spw_link_command_txdivcnt_o -> SpaceWire_Channel_B:spw_link_command_txdivcnt_i
	wire    [5:0] comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal;     // COMM_Pedreiro_v1_01_2:spw_timecode_tx_time_in_o -> SpaceWire_Channel_B:spw_timecode_tx_time_in_i
	wire          spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal;        // SpaceWire_Channel_B:spw_data_rx_status_rxflag_o -> COMM_Pedreiro_v1_01_2:spw_data_rx_status_rxflag_i
	wire    [1:0] comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal;     // COMM_Pedreiro_v1_01_2:spw_timecode_tx_ctrl_in_o -> SpaceWire_Channel_B:spw_timecode_tx_ctrl_in_i
	wire          comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_link_command_autostart_signal;  // COMM_Pedreiro_v1_01_2:spw_link_command_autostart_o -> SpaceWire_Channel_B:spw_link_command_autostart_i
	wire          spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errcred_signal;           // SpaceWire_Channel_B:spw_link_error_errcred_o -> COMM_Pedreiro_v1_01_2:spw_link_error_errcred_i
	wire          spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal;       // SpaceWire_Channel_D:spw_data_rx_status_rxvalid_o -> COMM_Pedreiro_v1_01_4:spw_data_rx_status_rxvalid_i
	wire    [7:0] comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal;  // COMM_Pedreiro_v1_01_4:spw_data_tx_command_txdata_o -> SpaceWire_Channel_D:spw_data_tx_command_txdata_i
	wire          spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errdisc_signal;           // SpaceWire_Channel_D:spw_link_error_errdisc_o -> COMM_Pedreiro_v1_01_4:spw_link_error_errdisc_i
	wire          spacewire_channel_d_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal;       // SpaceWire_Channel_D:spw_data_tx_status_txhalff_o -> COMM_Pedreiro_v1_01_4:spw_data_tx_status_txhalff_i
	wire          comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal; // COMM_Pedreiro_v1_01_4:spw_data_tx_command_txwrite_o -> SpaceWire_Channel_D:spw_data_tx_command_txwrite_i
	wire          spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal;         // SpaceWire_Channel_D:spw_timecode_rx_tick_out_o -> COMM_Pedreiro_v1_01_4:spw_timecode_rx_tick_out_i
	wire          spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal;       // SpaceWire_Channel_D:spw_data_rx_status_rxhalff_o -> COMM_Pedreiro_v1_01_4:spw_data_rx_status_rxhalff_i
	wire    [5:0] spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal;         // SpaceWire_Channel_D:spw_timecode_rx_time_out_o -> COMM_Pedreiro_v1_01_4:spw_timecode_rx_time_out_i
	wire          spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_connecting_signal;       // SpaceWire_Channel_D:spw_link_status_connecting_o -> COMM_Pedreiro_v1_01_4:spw_link_status_connecting_i
	wire    [7:0] spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal;        // SpaceWire_Channel_D:spw_data_rx_status_rxdata_o -> COMM_Pedreiro_v1_01_4:spw_data_rx_status_rxdata_i
	wire    [1:0] spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal;         // SpaceWire_Channel_D:spw_timecode_rx_ctrl_out_o -> COMM_Pedreiro_v1_01_4:spw_timecode_rx_ctrl_out_i
	wire          comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal;  // COMM_Pedreiro_v1_01_4:spw_data_tx_command_txflag_o -> SpaceWire_Channel_D:spw_data_tx_command_txflag_i
	wire          comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_link_command_linkstart_signal;  // COMM_Pedreiro_v1_01_4:spw_link_command_linkstart_o -> SpaceWire_Channel_D:spw_link_command_linkstart_i
	wire          comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal;  // COMM_Pedreiro_v1_01_4:spw_data_rx_command_rxread_o -> SpaceWire_Channel_D:spw_data_rx_command_rxread_i
	wire          spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_running_signal;          // SpaceWire_Channel_D:spw_link_status_running_o -> COMM_Pedreiro_v1_01_4:spw_link_status_running_i
	wire          spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_started_signal;          // SpaceWire_Channel_D:spw_link_status_started_o -> COMM_Pedreiro_v1_01_4:spw_link_status_started_i
	wire          spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errpar_signal;            // SpaceWire_Channel_D:spw_link_error_errpar_o -> COMM_Pedreiro_v1_01_4:spw_link_error_errpar_i
	wire          comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_link_command_linkdis_signal;    // COMM_Pedreiro_v1_01_4:spw_link_command_linkdis_o -> SpaceWire_Channel_D:spw_link_command_linkdis_i
	wire          spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_erresc_signal;            // SpaceWire_Channel_D:spw_link_error_erresc_o -> COMM_Pedreiro_v1_01_4:spw_link_error_erresc_i
	wire          spacewire_channel_d_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal;         // SpaceWire_Channel_D:spw_data_tx_status_txrdy_o -> COMM_Pedreiro_v1_01_4:spw_data_tx_status_txrdy_i
	wire          comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal;     // COMM_Pedreiro_v1_01_4:spw_timecode_tx_tick_in_o -> SpaceWire_Channel_D:spw_timecode_tx_tick_in_i
	wire    [7:0] comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal;   // COMM_Pedreiro_v1_01_4:spw_link_command_txdivcnt_o -> SpaceWire_Channel_D:spw_link_command_txdivcnt_i
	wire    [5:0] comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal;     // COMM_Pedreiro_v1_01_4:spw_timecode_tx_time_in_o -> SpaceWire_Channel_D:spw_timecode_tx_time_in_i
	wire          spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal;        // SpaceWire_Channel_D:spw_data_rx_status_rxflag_o -> COMM_Pedreiro_v1_01_4:spw_data_rx_status_rxflag_i
	wire    [1:0] comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal;     // COMM_Pedreiro_v1_01_4:spw_timecode_tx_ctrl_in_o -> SpaceWire_Channel_D:spw_timecode_tx_ctrl_in_i
	wire          comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_link_command_autostart_signal;  // COMM_Pedreiro_v1_01_4:spw_link_command_autostart_o -> SpaceWire_Channel_D:spw_link_command_autostart_i
	wire          spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errcred_signal;           // SpaceWire_Channel_D:spw_link_error_errcred_o -> COMM_Pedreiro_v1_01_4:spw_link_error_errcred_i
	wire          spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal;       // SpaceWire_Channel_F:spw_data_rx_status_rxvalid_o -> COMM_Pedreiro_v1_01_6:spw_data_rx_status_rxvalid_i
	wire    [7:0] comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal;  // COMM_Pedreiro_v1_01_6:spw_data_tx_command_txdata_o -> SpaceWire_Channel_F:spw_data_tx_command_txdata_i
	wire          spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errdisc_signal;           // SpaceWire_Channel_F:spw_link_error_errdisc_o -> COMM_Pedreiro_v1_01_6:spw_link_error_errdisc_i
	wire          spacewire_channel_f_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal;       // SpaceWire_Channel_F:spw_data_tx_status_txhalff_o -> COMM_Pedreiro_v1_01_6:spw_data_tx_status_txhalff_i
	wire          comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal; // COMM_Pedreiro_v1_01_6:spw_data_tx_command_txwrite_o -> SpaceWire_Channel_F:spw_data_tx_command_txwrite_i
	wire          spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal;         // SpaceWire_Channel_F:spw_timecode_rx_tick_out_o -> COMM_Pedreiro_v1_01_6:spw_timecode_rx_tick_out_i
	wire          spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal;       // SpaceWire_Channel_F:spw_data_rx_status_rxhalff_o -> COMM_Pedreiro_v1_01_6:spw_data_rx_status_rxhalff_i
	wire    [5:0] spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal;         // SpaceWire_Channel_F:spw_timecode_rx_time_out_o -> COMM_Pedreiro_v1_01_6:spw_timecode_rx_time_out_i
	wire          spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_connecting_signal;       // SpaceWire_Channel_F:spw_link_status_connecting_o -> COMM_Pedreiro_v1_01_6:spw_link_status_connecting_i
	wire    [7:0] spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal;        // SpaceWire_Channel_F:spw_data_rx_status_rxdata_o -> COMM_Pedreiro_v1_01_6:spw_data_rx_status_rxdata_i
	wire    [1:0] spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal;         // SpaceWire_Channel_F:spw_timecode_rx_ctrl_out_o -> COMM_Pedreiro_v1_01_6:spw_timecode_rx_ctrl_out_i
	wire          comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal;  // COMM_Pedreiro_v1_01_6:spw_data_tx_command_txflag_o -> SpaceWire_Channel_F:spw_data_tx_command_txflag_i
	wire          comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_link_command_linkstart_signal;  // COMM_Pedreiro_v1_01_6:spw_link_command_linkstart_o -> SpaceWire_Channel_F:spw_link_command_linkstart_i
	wire          comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal;  // COMM_Pedreiro_v1_01_6:spw_data_rx_command_rxread_o -> SpaceWire_Channel_F:spw_data_rx_command_rxread_i
	wire          spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_running_signal;          // SpaceWire_Channel_F:spw_link_status_running_o -> COMM_Pedreiro_v1_01_6:spw_link_status_running_i
	wire          spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_started_signal;          // SpaceWire_Channel_F:spw_link_status_started_o -> COMM_Pedreiro_v1_01_6:spw_link_status_started_i
	wire          spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errpar_signal;            // SpaceWire_Channel_F:spw_link_error_errpar_o -> COMM_Pedreiro_v1_01_6:spw_link_error_errpar_i
	wire          comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_link_command_linkdis_signal;    // COMM_Pedreiro_v1_01_6:spw_link_command_linkdis_o -> SpaceWire_Channel_F:spw_link_command_linkdis_i
	wire          spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_erresc_signal;            // SpaceWire_Channel_F:spw_link_error_erresc_o -> COMM_Pedreiro_v1_01_6:spw_link_error_erresc_i
	wire          spacewire_channel_f_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal;         // SpaceWire_Channel_F:spw_data_tx_status_txrdy_o -> COMM_Pedreiro_v1_01_6:spw_data_tx_status_txrdy_i
	wire          comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal;     // COMM_Pedreiro_v1_01_6:spw_timecode_tx_tick_in_o -> SpaceWire_Channel_F:spw_timecode_tx_tick_in_i
	wire    [7:0] comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal;   // COMM_Pedreiro_v1_01_6:spw_link_command_txdivcnt_o -> SpaceWire_Channel_F:spw_link_command_txdivcnt_i
	wire    [5:0] comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal;     // COMM_Pedreiro_v1_01_6:spw_timecode_tx_time_in_o -> SpaceWire_Channel_F:spw_timecode_tx_time_in_i
	wire          spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal;        // SpaceWire_Channel_F:spw_data_rx_status_rxflag_o -> COMM_Pedreiro_v1_01_6:spw_data_rx_status_rxflag_i
	wire    [1:0] comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal;     // COMM_Pedreiro_v1_01_6:spw_timecode_tx_ctrl_in_o -> SpaceWire_Channel_F:spw_timecode_tx_ctrl_in_i
	wire          comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_link_command_autostart_signal;  // COMM_Pedreiro_v1_01_6:spw_link_command_autostart_o -> SpaceWire_Channel_F:spw_link_command_autostart_i
	wire          spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errcred_signal;           // SpaceWire_Channel_F:spw_link_error_errcred_o -> COMM_Pedreiro_v1_01_6:spw_link_error_errcred_i
	wire          spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal;       // SpaceWire_Channel_C:spw_data_rx_status_rxvalid_o -> COMM_Pedreiro_v1_01_3:spw_data_rx_status_rxvalid_i
	wire    [7:0] comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal;  // COMM_Pedreiro_v1_01_3:spw_data_tx_command_txdata_o -> SpaceWire_Channel_C:spw_data_tx_command_txdata_i
	wire          spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errdisc_signal;           // SpaceWire_Channel_C:spw_link_error_errdisc_o -> COMM_Pedreiro_v1_01_3:spw_link_error_errdisc_i
	wire          spacewire_channel_c_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal;       // SpaceWire_Channel_C:spw_data_tx_status_txhalff_o -> COMM_Pedreiro_v1_01_3:spw_data_tx_status_txhalff_i
	wire          spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal;         // SpaceWire_Channel_C:spw_timecode_rx_tick_out_o -> COMM_Pedreiro_v1_01_3:spw_timecode_rx_tick_out_i
	wire          spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal;       // SpaceWire_Channel_C:spw_data_rx_status_rxhalff_o -> COMM_Pedreiro_v1_01_3:spw_data_rx_status_rxhalff_i
	wire          comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal; // COMM_Pedreiro_v1_01_3:spw_data_tx_command_txwrite_o -> SpaceWire_Channel_C:spw_data_tx_command_txwrite_i
	wire    [5:0] spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal;         // SpaceWire_Channel_C:spw_timecode_rx_time_out_o -> COMM_Pedreiro_v1_01_3:spw_timecode_rx_time_out_i
	wire          spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_connecting_signal;       // SpaceWire_Channel_C:spw_link_status_connecting_o -> COMM_Pedreiro_v1_01_3:spw_link_status_connecting_i
	wire    [7:0] spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal;        // SpaceWire_Channel_C:spw_data_rx_status_rxdata_o -> COMM_Pedreiro_v1_01_3:spw_data_rx_status_rxdata_i
	wire    [1:0] spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal;         // SpaceWire_Channel_C:spw_timecode_rx_ctrl_out_o -> COMM_Pedreiro_v1_01_3:spw_timecode_rx_ctrl_out_i
	wire          comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal;  // COMM_Pedreiro_v1_01_3:spw_data_tx_command_txflag_o -> SpaceWire_Channel_C:spw_data_tx_command_txflag_i
	wire          comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_link_command_linkstart_signal;  // COMM_Pedreiro_v1_01_3:spw_link_command_linkstart_o -> SpaceWire_Channel_C:spw_link_command_linkstart_i
	wire          comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal;  // COMM_Pedreiro_v1_01_3:spw_data_rx_command_rxread_o -> SpaceWire_Channel_C:spw_data_rx_command_rxread_i
	wire          spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_running_signal;          // SpaceWire_Channel_C:spw_link_status_running_o -> COMM_Pedreiro_v1_01_3:spw_link_status_running_i
	wire          spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_started_signal;          // SpaceWire_Channel_C:spw_link_status_started_o -> COMM_Pedreiro_v1_01_3:spw_link_status_started_i
	wire          spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errpar_signal;            // SpaceWire_Channel_C:spw_link_error_errpar_o -> COMM_Pedreiro_v1_01_3:spw_link_error_errpar_i
	wire          comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_link_command_linkdis_signal;    // COMM_Pedreiro_v1_01_3:spw_link_command_linkdis_o -> SpaceWire_Channel_C:spw_link_command_linkdis_i
	wire          spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_erresc_signal;            // SpaceWire_Channel_C:spw_link_error_erresc_o -> COMM_Pedreiro_v1_01_3:spw_link_error_erresc_i
	wire          spacewire_channel_c_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal;         // SpaceWire_Channel_C:spw_data_tx_status_txrdy_o -> COMM_Pedreiro_v1_01_3:spw_data_tx_status_txrdy_i
	wire          comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal;     // COMM_Pedreiro_v1_01_3:spw_timecode_tx_tick_in_o -> SpaceWire_Channel_C:spw_timecode_tx_tick_in_i
	wire    [7:0] comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal;   // COMM_Pedreiro_v1_01_3:spw_link_command_txdivcnt_o -> SpaceWire_Channel_C:spw_link_command_txdivcnt_i
	wire          spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal;        // SpaceWire_Channel_C:spw_data_rx_status_rxflag_o -> COMM_Pedreiro_v1_01_3:spw_data_rx_status_rxflag_i
	wire    [5:0] comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal;     // COMM_Pedreiro_v1_01_3:spw_timecode_tx_time_in_o -> SpaceWire_Channel_C:spw_timecode_tx_time_in_i
	wire    [1:0] comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal;     // COMM_Pedreiro_v1_01_3:spw_timecode_tx_ctrl_in_o -> SpaceWire_Channel_C:spw_timecode_tx_ctrl_in_i
	wire          comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_link_command_autostart_signal;  // COMM_Pedreiro_v1_01_3:spw_link_command_autostart_o -> SpaceWire_Channel_C:spw_link_command_autostart_i
	wire          spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errcred_signal;           // SpaceWire_Channel_C:spw_link_error_errcred_o -> COMM_Pedreiro_v1_01_3:spw_link_error_errcred_i
	wire          spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal;       // SpaceWire_Channel_E:spw_data_rx_status_rxvalid_o -> COMM_Pedreiro_v1_01_5:spw_data_rx_status_rxvalid_i
	wire    [7:0] comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal;  // COMM_Pedreiro_v1_01_5:spw_data_tx_command_txdata_o -> SpaceWire_Channel_E:spw_data_tx_command_txdata_i
	wire          spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errdisc_signal;           // SpaceWire_Channel_E:spw_link_error_errdisc_o -> COMM_Pedreiro_v1_01_5:spw_link_error_errdisc_i
	wire          spacewire_channel_e_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal;       // SpaceWire_Channel_E:spw_data_tx_status_txhalff_o -> COMM_Pedreiro_v1_01_5:spw_data_tx_status_txhalff_i
	wire          spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal;         // SpaceWire_Channel_E:spw_timecode_rx_tick_out_o -> COMM_Pedreiro_v1_01_5:spw_timecode_rx_tick_out_i
	wire          spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal;       // SpaceWire_Channel_E:spw_data_rx_status_rxhalff_o -> COMM_Pedreiro_v1_01_5:spw_data_rx_status_rxhalff_i
	wire          comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal; // COMM_Pedreiro_v1_01_5:spw_data_tx_command_txwrite_o -> SpaceWire_Channel_E:spw_data_tx_command_txwrite_i
	wire    [5:0] spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal;         // SpaceWire_Channel_E:spw_timecode_rx_time_out_o -> COMM_Pedreiro_v1_01_5:spw_timecode_rx_time_out_i
	wire          spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_connecting_signal;       // SpaceWire_Channel_E:spw_link_status_connecting_o -> COMM_Pedreiro_v1_01_5:spw_link_status_connecting_i
	wire    [7:0] spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal;        // SpaceWire_Channel_E:spw_data_rx_status_rxdata_o -> COMM_Pedreiro_v1_01_5:spw_data_rx_status_rxdata_i
	wire    [1:0] spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal;         // SpaceWire_Channel_E:spw_timecode_rx_ctrl_out_o -> COMM_Pedreiro_v1_01_5:spw_timecode_rx_ctrl_out_i
	wire          comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal;  // COMM_Pedreiro_v1_01_5:spw_data_tx_command_txflag_o -> SpaceWire_Channel_E:spw_data_tx_command_txflag_i
	wire          comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_link_command_linkstart_signal;  // COMM_Pedreiro_v1_01_5:spw_link_command_linkstart_o -> SpaceWire_Channel_E:spw_link_command_linkstart_i
	wire          comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal;  // COMM_Pedreiro_v1_01_5:spw_data_rx_command_rxread_o -> SpaceWire_Channel_E:spw_data_rx_command_rxread_i
	wire          spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_running_signal;          // SpaceWire_Channel_E:spw_link_status_running_o -> COMM_Pedreiro_v1_01_5:spw_link_status_running_i
	wire          spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_started_signal;          // SpaceWire_Channel_E:spw_link_status_started_o -> COMM_Pedreiro_v1_01_5:spw_link_status_started_i
	wire          spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errpar_signal;            // SpaceWire_Channel_E:spw_link_error_errpar_o -> COMM_Pedreiro_v1_01_5:spw_link_error_errpar_i
	wire          comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_link_command_linkdis_signal;    // COMM_Pedreiro_v1_01_5:spw_link_command_linkdis_o -> SpaceWire_Channel_E:spw_link_command_linkdis_i
	wire          spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_erresc_signal;            // SpaceWire_Channel_E:spw_link_error_erresc_o -> COMM_Pedreiro_v1_01_5:spw_link_error_erresc_i
	wire          spacewire_channel_e_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal;         // SpaceWire_Channel_E:spw_data_tx_status_txrdy_o -> COMM_Pedreiro_v1_01_5:spw_data_tx_status_txrdy_i
	wire          comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal;     // COMM_Pedreiro_v1_01_5:spw_timecode_tx_tick_in_o -> SpaceWire_Channel_E:spw_timecode_tx_tick_in_i
	wire    [7:0] comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal;   // COMM_Pedreiro_v1_01_5:spw_link_command_txdivcnt_o -> SpaceWire_Channel_E:spw_link_command_txdivcnt_i
	wire          spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal;        // SpaceWire_Channel_E:spw_data_rx_status_rxflag_o -> COMM_Pedreiro_v1_01_5:spw_data_rx_status_rxflag_i
	wire    [5:0] comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal;     // COMM_Pedreiro_v1_01_5:spw_timecode_tx_time_in_o -> SpaceWire_Channel_E:spw_timecode_tx_time_in_i
	wire    [1:0] comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal;     // COMM_Pedreiro_v1_01_5:spw_timecode_tx_ctrl_in_o -> SpaceWire_Channel_E:spw_timecode_tx_ctrl_in_i
	wire          comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_link_command_autostart_signal;  // COMM_Pedreiro_v1_01_5:spw_link_command_autostart_o -> SpaceWire_Channel_E:spw_link_command_autostart_i
	wire          spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errcred_signal;           // SpaceWire_Channel_E:spw_link_error_errcred_o -> COMM_Pedreiro_v1_01_5:spw_link_error_errcred_i
	wire          spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal;       // SpaceWire_Channel_G:spw_data_rx_status_rxvalid_o -> SpaceWire_Glutton_0:spw_data_rx_status_rxvalid_i
	wire    [7:0] spacewire_glutton_0_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal;    // SpaceWire_Glutton_0:spw_data_tx_command_txdata_o -> SpaceWire_Channel_G:spw_data_tx_command_txdata_i
	wire          spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errdisc_signal;           // SpaceWire_Channel_G:spw_link_error_errdisc_o -> SpaceWire_Glutton_0:spw_link_error_errdisc_i
	wire          spacewire_channel_g_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal;       // SpaceWire_Channel_G:spw_data_tx_status_txhalff_o -> SpaceWire_Glutton_0:spw_data_tx_status_txhalff_i
	wire          spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal;         // SpaceWire_Channel_G:spw_timecode_rx_tick_out_o -> SpaceWire_Glutton_0:spw_timecode_rx_tick_out_i
	wire          spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal;       // SpaceWire_Channel_G:spw_data_rx_status_rxhalff_o -> SpaceWire_Glutton_0:spw_data_rx_status_rxhalff_i
	wire          spacewire_glutton_0_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal;   // SpaceWire_Glutton_0:spw_data_tx_command_txwrite_o -> SpaceWire_Channel_G:spw_data_tx_command_txwrite_i
	wire    [5:0] spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal;         // SpaceWire_Channel_G:spw_timecode_rx_time_out_o -> SpaceWire_Glutton_0:spw_timecode_rx_time_out_i
	wire          spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_connecting_signal;       // SpaceWire_Channel_G:spw_link_status_connecting_o -> SpaceWire_Glutton_0:spw_link_status_connecting_i
	wire    [7:0] spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal;        // SpaceWire_Channel_G:spw_data_rx_status_rxdata_o -> SpaceWire_Glutton_0:spw_data_rx_status_rxdata_i
	wire    [1:0] spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal;         // SpaceWire_Channel_G:spw_timecode_rx_ctrl_out_o -> SpaceWire_Glutton_0:spw_timecode_rx_ctrl_out_i
	wire          spacewire_glutton_0_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal;    // SpaceWire_Glutton_0:spw_data_tx_command_txflag_o -> SpaceWire_Channel_G:spw_data_tx_command_txflag_i
	wire          spacewire_glutton_0_conduit_end_spacewire_controller_spw_link_command_linkstart_signal;    // SpaceWire_Glutton_0:spw_link_command_linkstart_o -> SpaceWire_Channel_G:spw_link_command_linkstart_i
	wire          spacewire_glutton_0_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal;    // SpaceWire_Glutton_0:spw_data_rx_command_rxread_o -> SpaceWire_Channel_G:spw_data_rx_command_rxread_i
	wire          spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_running_signal;          // SpaceWire_Channel_G:spw_link_status_running_o -> SpaceWire_Glutton_0:spw_link_status_running_i
	wire          spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_started_signal;          // SpaceWire_Channel_G:spw_link_status_started_o -> SpaceWire_Glutton_0:spw_link_status_started_i
	wire          spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errpar_signal;            // SpaceWire_Channel_G:spw_link_error_errpar_o -> SpaceWire_Glutton_0:spw_link_error_errpar_i
	wire          spacewire_glutton_0_conduit_end_spacewire_controller_spw_link_command_linkdis_signal;      // SpaceWire_Glutton_0:spw_link_command_linkdis_o -> SpaceWire_Channel_G:spw_link_command_linkdis_i
	wire          spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_erresc_signal;            // SpaceWire_Channel_G:spw_link_error_erresc_o -> SpaceWire_Glutton_0:spw_link_error_erresc_i
	wire          spacewire_channel_g_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal;         // SpaceWire_Channel_G:spw_data_tx_status_txrdy_o -> SpaceWire_Glutton_0:spw_data_tx_status_txrdy_i
	wire          spacewire_glutton_0_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal;       // SpaceWire_Glutton_0:spw_timecode_tx_tick_in_o -> SpaceWire_Channel_G:spw_timecode_tx_tick_in_i
	wire    [7:0] spacewire_glutton_0_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal;     // SpaceWire_Glutton_0:spw_link_command_txdivcnt_o -> SpaceWire_Channel_G:spw_link_command_txdivcnt_i
	wire          spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal;        // SpaceWire_Channel_G:spw_data_rx_status_rxflag_o -> SpaceWire_Glutton_0:spw_data_rx_status_rxflag_i
	wire    [5:0] spacewire_glutton_0_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal;       // SpaceWire_Glutton_0:spw_timecode_tx_time_in_o -> SpaceWire_Channel_G:spw_timecode_tx_time_in_i
	wire    [1:0] spacewire_glutton_0_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal;       // SpaceWire_Glutton_0:spw_timecode_tx_ctrl_in_o -> SpaceWire_Channel_G:spw_timecode_tx_ctrl_in_i
	wire          spacewire_glutton_0_conduit_end_spacewire_controller_spw_link_command_autostart_signal;    // SpaceWire_Glutton_0:spw_link_command_autostart_o -> SpaceWire_Channel_G:spw_link_command_autostart_i
	wire          spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errcred_signal;           // SpaceWire_Channel_G:spw_link_error_errcred_o -> SpaceWire_Glutton_0:spw_link_error_errcred_i
	wire          spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal;       // SpaceWire_Channel_H:spw_data_rx_status_rxvalid_o -> RMAP_Echoing_0:spw_data_rx_status_rxvalid_i
	wire    [7:0] rmap_echoing_0_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal;         // RMAP_Echoing_0:spw_data_tx_command_txdata_o -> SpaceWire_Channel_H:spw_data_tx_command_txdata_i
	wire          spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errdisc_signal;           // SpaceWire_Channel_H:spw_link_error_errdisc_o -> RMAP_Echoing_0:spw_link_error_errdisc_i
	wire          spacewire_channel_h_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal;       // SpaceWire_Channel_H:spw_data_tx_status_txhalff_o -> RMAP_Echoing_0:spw_data_tx_status_txhalff_i
	wire          spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal;         // SpaceWire_Channel_H:spw_timecode_rx_tick_out_o -> RMAP_Echoing_0:spw_timecode_rx_tick_out_i
	wire          spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal;       // SpaceWire_Channel_H:spw_data_rx_status_rxhalff_o -> RMAP_Echoing_0:spw_data_rx_status_rxhalff_i
	wire          rmap_echoing_0_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal;        // RMAP_Echoing_0:spw_data_tx_command_txwrite_o -> SpaceWire_Channel_H:spw_data_tx_command_txwrite_i
	wire    [5:0] spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal;         // SpaceWire_Channel_H:spw_timecode_rx_time_out_o -> RMAP_Echoing_0:spw_timecode_rx_time_out_i
	wire          spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_connecting_signal;       // SpaceWire_Channel_H:spw_link_status_connecting_o -> RMAP_Echoing_0:spw_link_status_connecting_i
	wire    [7:0] spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal;        // SpaceWire_Channel_H:spw_data_rx_status_rxdata_o -> RMAP_Echoing_0:spw_data_rx_status_rxdata_i
	wire    [1:0] spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal;         // SpaceWire_Channel_H:spw_timecode_rx_ctrl_out_o -> RMAP_Echoing_0:spw_timecode_rx_ctrl_out_i
	wire          rmap_echoing_0_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal;         // RMAP_Echoing_0:spw_data_tx_command_txflag_o -> SpaceWire_Channel_H:spw_data_tx_command_txflag_i
	wire          rmap_echoing_0_conduit_end_spacewire_controller_spw_link_command_linkstart_signal;         // RMAP_Echoing_0:spw_link_command_linkstart_o -> SpaceWire_Channel_H:spw_link_command_linkstart_i
	wire          rmap_echoing_0_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal;         // RMAP_Echoing_0:spw_data_rx_command_rxread_o -> SpaceWire_Channel_H:spw_data_rx_command_rxread_i
	wire          spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_running_signal;          // SpaceWire_Channel_H:spw_link_status_running_o -> RMAP_Echoing_0:spw_link_status_running_i
	wire          spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_started_signal;          // SpaceWire_Channel_H:spw_link_status_started_o -> RMAP_Echoing_0:spw_link_status_started_i
	wire          spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errpar_signal;            // SpaceWire_Channel_H:spw_link_error_errpar_o -> RMAP_Echoing_0:spw_link_error_errpar_i
	wire          rmap_echoing_0_conduit_end_spacewire_controller_spw_link_command_linkdis_signal;           // RMAP_Echoing_0:spw_link_command_linkdis_o -> SpaceWire_Channel_H:spw_link_command_linkdis_i
	wire          spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_erresc_signal;            // SpaceWire_Channel_H:spw_link_error_erresc_o -> RMAP_Echoing_0:spw_link_error_erresc_i
	wire          spacewire_channel_h_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal;         // SpaceWire_Channel_H:spw_data_tx_status_txrdy_o -> RMAP_Echoing_0:spw_data_tx_status_txrdy_i
	wire          rmap_echoing_0_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal;            // RMAP_Echoing_0:spw_timecode_tx_tick_in_o -> SpaceWire_Channel_H:spw_timecode_tx_tick_in_i
	wire    [7:0] rmap_echoing_0_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal;          // RMAP_Echoing_0:spw_link_command_txdivcnt_o -> SpaceWire_Channel_H:spw_link_command_txdivcnt_i
	wire          spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal;        // SpaceWire_Channel_H:spw_data_rx_status_rxflag_o -> RMAP_Echoing_0:spw_data_rx_status_rxflag_i
	wire    [5:0] rmap_echoing_0_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal;            // RMAP_Echoing_0:spw_timecode_tx_time_in_o -> SpaceWire_Channel_H:spw_timecode_tx_time_in_i
	wire    [1:0] rmap_echoing_0_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal;            // RMAP_Echoing_0:spw_timecode_tx_ctrl_in_o -> SpaceWire_Channel_H:spw_timecode_tx_ctrl_in_i
	wire          rmap_echoing_0_conduit_end_spacewire_controller_spw_link_command_autostart_signal;         // RMAP_Echoing_0:spw_link_command_autostart_o -> SpaceWire_Channel_H:spw_link_command_autostart_i
	wire          spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errcred_signal;           // SpaceWire_Channel_H:spw_link_error_errcred_o -> RMAP_Echoing_0:spw_link_error_errcred_i
	wire          ext_flash_tcm_data_outen;                                                                  // ext_flash:tcm_data_outen -> tristate_conduit_bridge_0:tcs_tcm_data_outen
	wire          ext_flash_tcm_request;                                                                     // ext_flash:tcm_request -> tristate_conduit_bridge_0:request
	wire          ext_flash_tcm_write_n_out;                                                                 // ext_flash:tcm_write_n_out -> tristate_conduit_bridge_0:tcs_tcm_write_n_out
	wire          ext_flash_tcm_read_n_out;                                                                  // ext_flash:tcm_read_n_out -> tristate_conduit_bridge_0:tcs_tcm_read_n_out
	wire          ext_flash_tcm_grant;                                                                       // tristate_conduit_bridge_0:grant -> ext_flash:tcm_grant
	wire          ext_flash_tcm_chipselect_n_out;                                                            // ext_flash:tcm_chipselect_n_out -> tristate_conduit_bridge_0:tcs_tcm_chipselect_n_out
	wire   [25:0] ext_flash_tcm_address_out;                                                                 // ext_flash:tcm_address_out -> tristate_conduit_bridge_0:tcs_tcm_address_out
	wire   [15:0] ext_flash_tcm_data_out;                                                                    // ext_flash:tcm_data_out -> tristate_conduit_bridge_0:tcs_tcm_data_out
	wire   [15:0] ext_flash_tcm_data_in;                                                                     // tristate_conduit_bridge_0:tcs_tcm_data_in -> ext_flash:tcm_data_in
	wire  [255:0] ftdi_usb3_0_avalon_master_data_readdata;                                                   // mm_interconnect_0:FTDI_USB3_0_avalon_master_data_readdata -> FTDI_USB3_0:avalon_master_data_readdata
	wire          ftdi_usb3_0_avalon_master_data_waitrequest;                                                // mm_interconnect_0:FTDI_USB3_0_avalon_master_data_waitrequest -> FTDI_USB3_0:avalon_master_data_waitrequest
	wire   [63:0] ftdi_usb3_0_avalon_master_data_address;                                                    // FTDI_USB3_0:avalon_master_data_address -> mm_interconnect_0:FTDI_USB3_0_avalon_master_data_address
	wire          ftdi_usb3_0_avalon_master_data_read;                                                       // FTDI_USB3_0:avalon_master_data_read -> mm_interconnect_0:FTDI_USB3_0_avalon_master_data_read
	wire          ftdi_usb3_0_avalon_master_data_write;                                                      // FTDI_USB3_0:avalon_master_data_write -> mm_interconnect_0:FTDI_USB3_0_avalon_master_data_write
	wire  [255:0] ftdi_usb3_0_avalon_master_data_writedata;                                                  // FTDI_USB3_0:avalon_master_data_writedata -> mm_interconnect_0:FTDI_USB3_0_avalon_master_data_writedata
	wire  [255:0] comm_pedreiro_v1_01_1_avalon_mm_left_buffer_master_readdata;                               // mm_interconnect_0:COMM_Pedreiro_v1_01_1_avalon_mm_left_buffer_master_readdata -> COMM_Pedreiro_v1_01_1:avm_left_buffer_readdata_i
	wire          comm_pedreiro_v1_01_1_avalon_mm_left_buffer_master_waitrequest;                            // mm_interconnect_0:COMM_Pedreiro_v1_01_1_avalon_mm_left_buffer_master_waitrequest -> COMM_Pedreiro_v1_01_1:avm_left_buffer_waitrequest_i
	wire   [63:0] comm_pedreiro_v1_01_1_avalon_mm_left_buffer_master_address;                                // COMM_Pedreiro_v1_01_1:avm_left_buffer_address_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_1_avalon_mm_left_buffer_master_address
	wire          comm_pedreiro_v1_01_1_avalon_mm_left_buffer_master_read;                                   // COMM_Pedreiro_v1_01_1:avm_left_buffer_read_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_1_avalon_mm_left_buffer_master_read
	wire  [255:0] comm_pedreiro_v1_01_2_avalon_mm_left_buffer_master_readdata;                               // mm_interconnect_0:COMM_Pedreiro_v1_01_2_avalon_mm_left_buffer_master_readdata -> COMM_Pedreiro_v1_01_2:avm_left_buffer_readdata_i
	wire          comm_pedreiro_v1_01_2_avalon_mm_left_buffer_master_waitrequest;                            // mm_interconnect_0:COMM_Pedreiro_v1_01_2_avalon_mm_left_buffer_master_waitrequest -> COMM_Pedreiro_v1_01_2:avm_left_buffer_waitrequest_i
	wire   [63:0] comm_pedreiro_v1_01_2_avalon_mm_left_buffer_master_address;                                // COMM_Pedreiro_v1_01_2:avm_left_buffer_address_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_2_avalon_mm_left_buffer_master_address
	wire          comm_pedreiro_v1_01_2_avalon_mm_left_buffer_master_read;                                   // COMM_Pedreiro_v1_01_2:avm_left_buffer_read_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_2_avalon_mm_left_buffer_master_read
	wire  [255:0] comm_pedreiro_v1_01_3_avalon_mm_left_buffer_master_readdata;                               // mm_interconnect_0:COMM_Pedreiro_v1_01_3_avalon_mm_left_buffer_master_readdata -> COMM_Pedreiro_v1_01_3:avm_left_buffer_readdata_i
	wire          comm_pedreiro_v1_01_3_avalon_mm_left_buffer_master_waitrequest;                            // mm_interconnect_0:COMM_Pedreiro_v1_01_3_avalon_mm_left_buffer_master_waitrequest -> COMM_Pedreiro_v1_01_3:avm_left_buffer_waitrequest_i
	wire   [63:0] comm_pedreiro_v1_01_3_avalon_mm_left_buffer_master_address;                                // COMM_Pedreiro_v1_01_3:avm_left_buffer_address_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_3_avalon_mm_left_buffer_master_address
	wire          comm_pedreiro_v1_01_3_avalon_mm_left_buffer_master_read;                                   // COMM_Pedreiro_v1_01_3:avm_left_buffer_read_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_3_avalon_mm_left_buffer_master_read
	wire  [255:0] comm_pedreiro_v1_01_4_avalon_mm_left_buffer_master_readdata;                               // mm_interconnect_0:COMM_Pedreiro_v1_01_4_avalon_mm_left_buffer_master_readdata -> COMM_Pedreiro_v1_01_4:avm_left_buffer_readdata_i
	wire          comm_pedreiro_v1_01_4_avalon_mm_left_buffer_master_waitrequest;                            // mm_interconnect_0:COMM_Pedreiro_v1_01_4_avalon_mm_left_buffer_master_waitrequest -> COMM_Pedreiro_v1_01_4:avm_left_buffer_waitrequest_i
	wire   [63:0] comm_pedreiro_v1_01_4_avalon_mm_left_buffer_master_address;                                // COMM_Pedreiro_v1_01_4:avm_left_buffer_address_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_4_avalon_mm_left_buffer_master_address
	wire          comm_pedreiro_v1_01_4_avalon_mm_left_buffer_master_read;                                   // COMM_Pedreiro_v1_01_4:avm_left_buffer_read_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_4_avalon_mm_left_buffer_master_read
	wire  [255:0] comm_pedreiro_v1_01_5_avalon_mm_left_buffer_master_readdata;                               // mm_interconnect_0:COMM_Pedreiro_v1_01_5_avalon_mm_left_buffer_master_readdata -> COMM_Pedreiro_v1_01_5:avm_left_buffer_readdata_i
	wire          comm_pedreiro_v1_01_5_avalon_mm_left_buffer_master_waitrequest;                            // mm_interconnect_0:COMM_Pedreiro_v1_01_5_avalon_mm_left_buffer_master_waitrequest -> COMM_Pedreiro_v1_01_5:avm_left_buffer_waitrequest_i
	wire   [63:0] comm_pedreiro_v1_01_5_avalon_mm_left_buffer_master_address;                                // COMM_Pedreiro_v1_01_5:avm_left_buffer_address_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_5_avalon_mm_left_buffer_master_address
	wire          comm_pedreiro_v1_01_5_avalon_mm_left_buffer_master_read;                                   // COMM_Pedreiro_v1_01_5:avm_left_buffer_read_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_5_avalon_mm_left_buffer_master_read
	wire  [255:0] comm_pedreiro_v1_01_6_avalon_mm_left_buffer_master_readdata;                               // mm_interconnect_0:COMM_Pedreiro_v1_01_6_avalon_mm_left_buffer_master_readdata -> COMM_Pedreiro_v1_01_6:avm_left_buffer_readdata_i
	wire          comm_pedreiro_v1_01_6_avalon_mm_left_buffer_master_waitrequest;                            // mm_interconnect_0:COMM_Pedreiro_v1_01_6_avalon_mm_left_buffer_master_waitrequest -> COMM_Pedreiro_v1_01_6:avm_left_buffer_waitrequest_i
	wire   [63:0] comm_pedreiro_v1_01_6_avalon_mm_left_buffer_master_address;                                // COMM_Pedreiro_v1_01_6:avm_left_buffer_address_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_6_avalon_mm_left_buffer_master_address
	wire          comm_pedreiro_v1_01_6_avalon_mm_left_buffer_master_read;                                   // COMM_Pedreiro_v1_01_6:avm_left_buffer_read_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_6_avalon_mm_left_buffer_master_read
	wire  [255:0] comm_pedreiro_v1_01_1_avalon_mm_right_buffer_master_readdata;                              // mm_interconnect_0:COMM_Pedreiro_v1_01_1_avalon_mm_right_buffer_master_readdata -> COMM_Pedreiro_v1_01_1:avm_right_buffer_readdata_i
	wire          comm_pedreiro_v1_01_1_avalon_mm_right_buffer_master_waitrequest;                           // mm_interconnect_0:COMM_Pedreiro_v1_01_1_avalon_mm_right_buffer_master_waitrequest -> COMM_Pedreiro_v1_01_1:avm_right_buffer_waitrequest_i
	wire   [63:0] comm_pedreiro_v1_01_1_avalon_mm_right_buffer_master_address;                               // COMM_Pedreiro_v1_01_1:avm_right_buffer_address_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_1_avalon_mm_right_buffer_master_address
	wire          comm_pedreiro_v1_01_1_avalon_mm_right_buffer_master_read;                                  // COMM_Pedreiro_v1_01_1:avm_right_buffer_read_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_1_avalon_mm_right_buffer_master_read
	wire  [255:0] comm_pedreiro_v1_01_2_avalon_mm_right_buffer_master_readdata;                              // mm_interconnect_0:COMM_Pedreiro_v1_01_2_avalon_mm_right_buffer_master_readdata -> COMM_Pedreiro_v1_01_2:avm_right_buffer_readdata_i
	wire          comm_pedreiro_v1_01_2_avalon_mm_right_buffer_master_waitrequest;                           // mm_interconnect_0:COMM_Pedreiro_v1_01_2_avalon_mm_right_buffer_master_waitrequest -> COMM_Pedreiro_v1_01_2:avm_right_buffer_waitrequest_i
	wire   [63:0] comm_pedreiro_v1_01_2_avalon_mm_right_buffer_master_address;                               // COMM_Pedreiro_v1_01_2:avm_right_buffer_address_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_2_avalon_mm_right_buffer_master_address
	wire          comm_pedreiro_v1_01_2_avalon_mm_right_buffer_master_read;                                  // COMM_Pedreiro_v1_01_2:avm_right_buffer_read_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_2_avalon_mm_right_buffer_master_read
	wire  [255:0] comm_pedreiro_v1_01_3_avalon_mm_right_buffer_master_readdata;                              // mm_interconnect_0:COMM_Pedreiro_v1_01_3_avalon_mm_right_buffer_master_readdata -> COMM_Pedreiro_v1_01_3:avm_right_buffer_readdata_i
	wire          comm_pedreiro_v1_01_3_avalon_mm_right_buffer_master_waitrequest;                           // mm_interconnect_0:COMM_Pedreiro_v1_01_3_avalon_mm_right_buffer_master_waitrequest -> COMM_Pedreiro_v1_01_3:avm_right_buffer_waitrequest_i
	wire   [63:0] comm_pedreiro_v1_01_3_avalon_mm_right_buffer_master_address;                               // COMM_Pedreiro_v1_01_3:avm_right_buffer_address_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_3_avalon_mm_right_buffer_master_address
	wire          comm_pedreiro_v1_01_3_avalon_mm_right_buffer_master_read;                                  // COMM_Pedreiro_v1_01_3:avm_right_buffer_read_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_3_avalon_mm_right_buffer_master_read
	wire  [255:0] comm_pedreiro_v1_01_4_avalon_mm_right_buffer_master_readdata;                              // mm_interconnect_0:COMM_Pedreiro_v1_01_4_avalon_mm_right_buffer_master_readdata -> COMM_Pedreiro_v1_01_4:avm_right_buffer_readdata_i
	wire          comm_pedreiro_v1_01_4_avalon_mm_right_buffer_master_waitrequest;                           // mm_interconnect_0:COMM_Pedreiro_v1_01_4_avalon_mm_right_buffer_master_waitrequest -> COMM_Pedreiro_v1_01_4:avm_right_buffer_waitrequest_i
	wire   [63:0] comm_pedreiro_v1_01_4_avalon_mm_right_buffer_master_address;                               // COMM_Pedreiro_v1_01_4:avm_right_buffer_address_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_4_avalon_mm_right_buffer_master_address
	wire          comm_pedreiro_v1_01_4_avalon_mm_right_buffer_master_read;                                  // COMM_Pedreiro_v1_01_4:avm_right_buffer_read_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_4_avalon_mm_right_buffer_master_read
	wire  [255:0] comm_pedreiro_v1_01_5_avalon_mm_right_buffer_master_readdata;                              // mm_interconnect_0:COMM_Pedreiro_v1_01_5_avalon_mm_right_buffer_master_readdata -> COMM_Pedreiro_v1_01_5:avm_right_buffer_readdata_i
	wire          comm_pedreiro_v1_01_5_avalon_mm_right_buffer_master_waitrequest;                           // mm_interconnect_0:COMM_Pedreiro_v1_01_5_avalon_mm_right_buffer_master_waitrequest -> COMM_Pedreiro_v1_01_5:avm_right_buffer_waitrequest_i
	wire   [63:0] comm_pedreiro_v1_01_5_avalon_mm_right_buffer_master_address;                               // COMM_Pedreiro_v1_01_5:avm_right_buffer_address_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_5_avalon_mm_right_buffer_master_address
	wire          comm_pedreiro_v1_01_5_avalon_mm_right_buffer_master_read;                                  // COMM_Pedreiro_v1_01_5:avm_right_buffer_read_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_5_avalon_mm_right_buffer_master_read
	wire  [255:0] comm_pedreiro_v1_01_6_avalon_mm_right_buffer_master_readdata;                              // mm_interconnect_0:COMM_Pedreiro_v1_01_6_avalon_mm_right_buffer_master_readdata -> COMM_Pedreiro_v1_01_6:avm_right_buffer_readdata_i
	wire          comm_pedreiro_v1_01_6_avalon_mm_right_buffer_master_waitrequest;                           // mm_interconnect_0:COMM_Pedreiro_v1_01_6_avalon_mm_right_buffer_master_waitrequest -> COMM_Pedreiro_v1_01_6:avm_right_buffer_waitrequest_i
	wire   [63:0] comm_pedreiro_v1_01_6_avalon_mm_right_buffer_master_address;                               // COMM_Pedreiro_v1_01_6:avm_right_buffer_address_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_6_avalon_mm_right_buffer_master_address
	wire          comm_pedreiro_v1_01_6_avalon_mm_right_buffer_master_read;                                  // COMM_Pedreiro_v1_01_6:avm_right_buffer_read_o -> mm_interconnect_0:COMM_Pedreiro_v1_01_6_avalon_mm_right_buffer_master_read
	wire    [7:0] rmap_mem_nfee_comm_1_avalon_mm_rmap_master_readdata;                                       // mm_interconnect_0:rmap_mem_nfee_comm_1_avalon_mm_rmap_master_readdata -> rmap_mem_nfee_comm_1:avm_rmap_readdata_i
	wire          rmap_mem_nfee_comm_1_avalon_mm_rmap_master_waitrequest;                                    // mm_interconnect_0:rmap_mem_nfee_comm_1_avalon_mm_rmap_master_waitrequest -> rmap_mem_nfee_comm_1:avm_rmap_waitrequest_i
	wire   [63:0] rmap_mem_nfee_comm_1_avalon_mm_rmap_master_address;                                        // rmap_mem_nfee_comm_1:avm_rmap_address_o -> mm_interconnect_0:rmap_mem_nfee_comm_1_avalon_mm_rmap_master_address
	wire          rmap_mem_nfee_comm_1_avalon_mm_rmap_master_read;                                           // rmap_mem_nfee_comm_1:avm_rmap_read_o -> mm_interconnect_0:rmap_mem_nfee_comm_1_avalon_mm_rmap_master_read
	wire          rmap_mem_nfee_comm_1_avalon_mm_rmap_master_write;                                          // rmap_mem_nfee_comm_1:avm_rmap_write_o -> mm_interconnect_0:rmap_mem_nfee_comm_1_avalon_mm_rmap_master_write
	wire    [7:0] rmap_mem_nfee_comm_1_avalon_mm_rmap_master_writedata;                                      // rmap_mem_nfee_comm_1:avm_rmap_writedata_o -> mm_interconnect_0:rmap_mem_nfee_comm_1_avalon_mm_rmap_master_writedata
	wire    [7:0] rmap_mem_nfee_comm_2_avalon_mm_rmap_master_readdata;                                       // mm_interconnect_0:rmap_mem_nfee_comm_2_avalon_mm_rmap_master_readdata -> rmap_mem_nfee_comm_2:avm_rmap_readdata_i
	wire          rmap_mem_nfee_comm_2_avalon_mm_rmap_master_waitrequest;                                    // mm_interconnect_0:rmap_mem_nfee_comm_2_avalon_mm_rmap_master_waitrequest -> rmap_mem_nfee_comm_2:avm_rmap_waitrequest_i
	wire   [63:0] rmap_mem_nfee_comm_2_avalon_mm_rmap_master_address;                                        // rmap_mem_nfee_comm_2:avm_rmap_address_o -> mm_interconnect_0:rmap_mem_nfee_comm_2_avalon_mm_rmap_master_address
	wire          rmap_mem_nfee_comm_2_avalon_mm_rmap_master_read;                                           // rmap_mem_nfee_comm_2:avm_rmap_read_o -> mm_interconnect_0:rmap_mem_nfee_comm_2_avalon_mm_rmap_master_read
	wire          rmap_mem_nfee_comm_2_avalon_mm_rmap_master_write;                                          // rmap_mem_nfee_comm_2:avm_rmap_write_o -> mm_interconnect_0:rmap_mem_nfee_comm_2_avalon_mm_rmap_master_write
	wire    [7:0] rmap_mem_nfee_comm_2_avalon_mm_rmap_master_writedata;                                      // rmap_mem_nfee_comm_2:avm_rmap_writedata_o -> mm_interconnect_0:rmap_mem_nfee_comm_2_avalon_mm_rmap_master_writedata
	wire    [7:0] rmap_mem_nfee_comm_3_avalon_mm_rmap_master_readdata;                                       // mm_interconnect_0:rmap_mem_nfee_comm_3_avalon_mm_rmap_master_readdata -> rmap_mem_nfee_comm_3:avm_rmap_readdata_i
	wire          rmap_mem_nfee_comm_3_avalon_mm_rmap_master_waitrequest;                                    // mm_interconnect_0:rmap_mem_nfee_comm_3_avalon_mm_rmap_master_waitrequest -> rmap_mem_nfee_comm_3:avm_rmap_waitrequest_i
	wire   [63:0] rmap_mem_nfee_comm_3_avalon_mm_rmap_master_address;                                        // rmap_mem_nfee_comm_3:avm_rmap_address_o -> mm_interconnect_0:rmap_mem_nfee_comm_3_avalon_mm_rmap_master_address
	wire          rmap_mem_nfee_comm_3_avalon_mm_rmap_master_read;                                           // rmap_mem_nfee_comm_3:avm_rmap_read_o -> mm_interconnect_0:rmap_mem_nfee_comm_3_avalon_mm_rmap_master_read
	wire          rmap_mem_nfee_comm_3_avalon_mm_rmap_master_write;                                          // rmap_mem_nfee_comm_3:avm_rmap_write_o -> mm_interconnect_0:rmap_mem_nfee_comm_3_avalon_mm_rmap_master_write
	wire    [7:0] rmap_mem_nfee_comm_3_avalon_mm_rmap_master_writedata;                                      // rmap_mem_nfee_comm_3:avm_rmap_writedata_o -> mm_interconnect_0:rmap_mem_nfee_comm_3_avalon_mm_rmap_master_writedata
	wire    [7:0] rmap_mem_nfee_comm_4_avalon_mm_rmap_master_readdata;                                       // mm_interconnect_0:rmap_mem_nfee_comm_4_avalon_mm_rmap_master_readdata -> rmap_mem_nfee_comm_4:avm_rmap_readdata_i
	wire          rmap_mem_nfee_comm_4_avalon_mm_rmap_master_waitrequest;                                    // mm_interconnect_0:rmap_mem_nfee_comm_4_avalon_mm_rmap_master_waitrequest -> rmap_mem_nfee_comm_4:avm_rmap_waitrequest_i
	wire   [63:0] rmap_mem_nfee_comm_4_avalon_mm_rmap_master_address;                                        // rmap_mem_nfee_comm_4:avm_rmap_address_o -> mm_interconnect_0:rmap_mem_nfee_comm_4_avalon_mm_rmap_master_address
	wire          rmap_mem_nfee_comm_4_avalon_mm_rmap_master_read;                                           // rmap_mem_nfee_comm_4:avm_rmap_read_o -> mm_interconnect_0:rmap_mem_nfee_comm_4_avalon_mm_rmap_master_read
	wire          rmap_mem_nfee_comm_4_avalon_mm_rmap_master_write;                                          // rmap_mem_nfee_comm_4:avm_rmap_write_o -> mm_interconnect_0:rmap_mem_nfee_comm_4_avalon_mm_rmap_master_write
	wire    [7:0] rmap_mem_nfee_comm_4_avalon_mm_rmap_master_writedata;                                      // rmap_mem_nfee_comm_4:avm_rmap_writedata_o -> mm_interconnect_0:rmap_mem_nfee_comm_4_avalon_mm_rmap_master_writedata
	wire    [7:0] rmap_mem_nfee_comm_5_avalon_mm_rmap_master_readdata;                                       // mm_interconnect_0:rmap_mem_nfee_comm_5_avalon_mm_rmap_master_readdata -> rmap_mem_nfee_comm_5:avm_rmap_readdata_i
	wire          rmap_mem_nfee_comm_5_avalon_mm_rmap_master_waitrequest;                                    // mm_interconnect_0:rmap_mem_nfee_comm_5_avalon_mm_rmap_master_waitrequest -> rmap_mem_nfee_comm_5:avm_rmap_waitrequest_i
	wire   [63:0] rmap_mem_nfee_comm_5_avalon_mm_rmap_master_address;                                        // rmap_mem_nfee_comm_5:avm_rmap_address_o -> mm_interconnect_0:rmap_mem_nfee_comm_5_avalon_mm_rmap_master_address
	wire          rmap_mem_nfee_comm_5_avalon_mm_rmap_master_read;                                           // rmap_mem_nfee_comm_5:avm_rmap_read_o -> mm_interconnect_0:rmap_mem_nfee_comm_5_avalon_mm_rmap_master_read
	wire          rmap_mem_nfee_comm_5_avalon_mm_rmap_master_write;                                          // rmap_mem_nfee_comm_5:avm_rmap_write_o -> mm_interconnect_0:rmap_mem_nfee_comm_5_avalon_mm_rmap_master_write
	wire    [7:0] rmap_mem_nfee_comm_5_avalon_mm_rmap_master_writedata;                                      // rmap_mem_nfee_comm_5:avm_rmap_writedata_o -> mm_interconnect_0:rmap_mem_nfee_comm_5_avalon_mm_rmap_master_writedata
	wire    [7:0] rmap_mem_nfee_comm_6_avalon_mm_rmap_master_readdata;                                       // mm_interconnect_0:rmap_mem_nfee_comm_6_avalon_mm_rmap_master_readdata -> rmap_mem_nfee_comm_6:avm_rmap_readdata_i
	wire          rmap_mem_nfee_comm_6_avalon_mm_rmap_master_waitrequest;                                    // mm_interconnect_0:rmap_mem_nfee_comm_6_avalon_mm_rmap_master_waitrequest -> rmap_mem_nfee_comm_6:avm_rmap_waitrequest_i
	wire   [63:0] rmap_mem_nfee_comm_6_avalon_mm_rmap_master_address;                                        // rmap_mem_nfee_comm_6:avm_rmap_address_o -> mm_interconnect_0:rmap_mem_nfee_comm_6_avalon_mm_rmap_master_address
	wire          rmap_mem_nfee_comm_6_avalon_mm_rmap_master_read;                                           // rmap_mem_nfee_comm_6:avm_rmap_read_o -> mm_interconnect_0:rmap_mem_nfee_comm_6_avalon_mm_rmap_master_read
	wire          rmap_mem_nfee_comm_6_avalon_mm_rmap_master_write;                                          // rmap_mem_nfee_comm_6:avm_rmap_write_o -> mm_interconnect_0:rmap_mem_nfee_comm_6_avalon_mm_rmap_master_write
	wire    [7:0] rmap_mem_nfee_comm_6_avalon_mm_rmap_master_writedata;                                      // rmap_mem_nfee_comm_6:avm_rmap_writedata_o -> mm_interconnect_0:rmap_mem_nfee_comm_6_avalon_mm_rmap_master_writedata
	wire          ddr2_address_span_extender_expanded_master_waitrequest;                                    // mm_interconnect_0:ddr2_address_span_extender_expanded_master_waitrequest -> ddr2_address_span_extender:avm_m0_waitrequest
	wire   [31:0] ddr2_address_span_extender_expanded_master_readdata;                                       // mm_interconnect_0:ddr2_address_span_extender_expanded_master_readdata -> ddr2_address_span_extender:avm_m0_readdata
	wire   [31:0] ddr2_address_span_extender_expanded_master_address;                                        // ddr2_address_span_extender:avm_m0_address -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_address
	wire          ddr2_address_span_extender_expanded_master_read;                                           // ddr2_address_span_extender:avm_m0_read -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_read
	wire    [3:0] ddr2_address_span_extender_expanded_master_byteenable;                                     // ddr2_address_span_extender:avm_m0_byteenable -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_byteenable
	wire          ddr2_address_span_extender_expanded_master_readdatavalid;                                  // mm_interconnect_0:ddr2_address_span_extender_expanded_master_readdatavalid -> ddr2_address_span_extender:avm_m0_readdatavalid
	wire          ddr2_address_span_extender_expanded_master_write;                                          // ddr2_address_span_extender:avm_m0_write -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_write
	wire   [31:0] ddr2_address_span_extender_expanded_master_writedata;                                      // ddr2_address_span_extender:avm_m0_writedata -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_writedata
	wire    [7:0] ddr2_address_span_extender_expanded_master_burstcount;                                     // ddr2_address_span_extender:avm_m0_burstcount -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_burstcount
	wire          mm_interconnect_0_m2_ddr2_memory_avl_beginbursttransfer;                                   // mm_interconnect_0:m2_ddr2_memory_avl_beginbursttransfer -> m2_ddr2_memory:avl_burstbegin
	wire  [255:0] mm_interconnect_0_m2_ddr2_memory_avl_readdata;                                             // m2_ddr2_memory:avl_rdata -> mm_interconnect_0:m2_ddr2_memory_avl_readdata
	wire          mm_interconnect_0_m2_ddr2_memory_avl_waitrequest;                                          // m2_ddr2_memory:avl_ready -> mm_interconnect_0:m2_ddr2_memory_avl_waitrequest
	wire   [25:0] mm_interconnect_0_m2_ddr2_memory_avl_address;                                              // mm_interconnect_0:m2_ddr2_memory_avl_address -> m2_ddr2_memory:avl_addr
	wire          mm_interconnect_0_m2_ddr2_memory_avl_read;                                                 // mm_interconnect_0:m2_ddr2_memory_avl_read -> m2_ddr2_memory:avl_read_req
	wire   [31:0] mm_interconnect_0_m2_ddr2_memory_avl_byteenable;                                           // mm_interconnect_0:m2_ddr2_memory_avl_byteenable -> m2_ddr2_memory:avl_be
	wire          mm_interconnect_0_m2_ddr2_memory_avl_readdatavalid;                                        // m2_ddr2_memory:avl_rdata_valid -> mm_interconnect_0:m2_ddr2_memory_avl_readdatavalid
	wire          mm_interconnect_0_m2_ddr2_memory_avl_write;                                                // mm_interconnect_0:m2_ddr2_memory_avl_write -> m2_ddr2_memory:avl_write_req
	wire  [255:0] mm_interconnect_0_m2_ddr2_memory_avl_writedata;                                            // mm_interconnect_0:m2_ddr2_memory_avl_writedata -> m2_ddr2_memory:avl_wdata
	wire    [7:0] mm_interconnect_0_m2_ddr2_memory_avl_burstcount;                                           // mm_interconnect_0:m2_ddr2_memory_avl_burstcount -> m2_ddr2_memory:avl_size
	wire  [255:0] mm_interconnect_0_m1_clock_bridge_s0_readdata;                                             // m1_clock_bridge:s0_readdata -> mm_interconnect_0:m1_clock_bridge_s0_readdata
	wire          mm_interconnect_0_m1_clock_bridge_s0_waitrequest;                                          // m1_clock_bridge:s0_waitrequest -> mm_interconnect_0:m1_clock_bridge_s0_waitrequest
	wire          mm_interconnect_0_m1_clock_bridge_s0_debugaccess;                                          // mm_interconnect_0:m1_clock_bridge_s0_debugaccess -> m1_clock_bridge:s0_debugaccess
	wire   [30:0] mm_interconnect_0_m1_clock_bridge_s0_address;                                              // mm_interconnect_0:m1_clock_bridge_s0_address -> m1_clock_bridge:s0_address
	wire          mm_interconnect_0_m1_clock_bridge_s0_read;                                                 // mm_interconnect_0:m1_clock_bridge_s0_read -> m1_clock_bridge:s0_read
	wire   [31:0] mm_interconnect_0_m1_clock_bridge_s0_byteenable;                                           // mm_interconnect_0:m1_clock_bridge_s0_byteenable -> m1_clock_bridge:s0_byteenable
	wire          mm_interconnect_0_m1_clock_bridge_s0_readdatavalid;                                        // m1_clock_bridge:s0_readdatavalid -> mm_interconnect_0:m1_clock_bridge_s0_readdatavalid
	wire          mm_interconnect_0_m1_clock_bridge_s0_write;                                                // mm_interconnect_0:m1_clock_bridge_s0_write -> m1_clock_bridge:s0_write
	wire  [255:0] mm_interconnect_0_m1_clock_bridge_s0_writedata;                                            // mm_interconnect_0:m1_clock_bridge_s0_writedata -> m1_clock_bridge:s0_writedata
	wire    [2:0] mm_interconnect_0_m1_clock_bridge_s0_burstcount;                                           // mm_interconnect_0:m1_clock_bridge_s0_burstcount -> m1_clock_bridge:s0_burstcount
	wire   [31:0] nios2_gen2_0_data_master_readdata;                                                         // mm_interconnect_1:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire          nios2_gen2_0_data_master_waitrequest;                                                      // mm_interconnect_1:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire          nios2_gen2_0_data_master_debugaccess;                                                      // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:nios2_gen2_0_data_master_debugaccess
	wire   [31:0] nios2_gen2_0_data_master_address;                                                          // nios2_gen2_0:d_address -> mm_interconnect_1:nios2_gen2_0_data_master_address
	wire    [3:0] nios2_gen2_0_data_master_byteenable;                                                       // nios2_gen2_0:d_byteenable -> mm_interconnect_1:nios2_gen2_0_data_master_byteenable
	wire          nios2_gen2_0_data_master_read;                                                             // nios2_gen2_0:d_read -> mm_interconnect_1:nios2_gen2_0_data_master_read
	wire          nios2_gen2_0_data_master_write;                                                            // nios2_gen2_0:d_write -> mm_interconnect_1:nios2_gen2_0_data_master_write
	wire   [31:0] nios2_gen2_0_data_master_writedata;                                                        // nios2_gen2_0:d_writedata -> mm_interconnect_1:nios2_gen2_0_data_master_writedata
	wire   [31:0] nios2_gen2_0_instruction_master_readdata;                                                  // mm_interconnect_1:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire          nios2_gen2_0_instruction_master_waitrequest;                                               // mm_interconnect_1:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire   [31:0] nios2_gen2_0_instruction_master_address;                                                   // nios2_gen2_0:i_address -> mm_interconnect_1:nios2_gen2_0_instruction_master_address
	wire          nios2_gen2_0_instruction_master_read;                                                      // nios2_gen2_0:i_read -> mm_interconnect_1:nios2_gen2_0_instruction_master_read
	wire          nios2_gen2_0_instruction_master_readdatavalid;                                             // mm_interconnect_1:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire    [3:0] nios2_gen2_0_instruction_master_burstcount;                                                // nios2_gen2_0:i_burstcount -> mm_interconnect_1:nios2_gen2_0_instruction_master_burstcount
	wire          mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect;                                // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire   [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata;                                  // jtag_uart_0:av_readdata -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_readdata
	wire          mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest;                               // jtag_uart_0:av_waitrequest -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address;                                   // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire          mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read;                                      // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire          mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write;                                     // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire   [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata;                                 // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [31:0] mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_readdata;                       // rmap_mem_nfee_comm_1:avs_0_rmap_readdata_o -> mm_interconnect_1:rmap_mem_nfee_comm_1_avalon_rmap_slave_0_readdata
	wire          mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_waitrequest;                    // rmap_mem_nfee_comm_1:avs_0_rmap_waitrequest_o -> mm_interconnect_1:rmap_mem_nfee_comm_1_avalon_rmap_slave_0_waitrequest
	wire   [11:0] mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_address;                        // mm_interconnect_1:rmap_mem_nfee_comm_1_avalon_rmap_slave_0_address -> rmap_mem_nfee_comm_1:avs_0_rmap_address_i
	wire          mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_read;                           // mm_interconnect_1:rmap_mem_nfee_comm_1_avalon_rmap_slave_0_read -> rmap_mem_nfee_comm_1:avs_0_rmap_read_i
	wire    [3:0] mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_byteenable;                     // mm_interconnect_1:rmap_mem_nfee_comm_1_avalon_rmap_slave_0_byteenable -> rmap_mem_nfee_comm_1:avs_0_rmap_byteenable_i
	wire          mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_write;                          // mm_interconnect_1:rmap_mem_nfee_comm_1_avalon_rmap_slave_0_write -> rmap_mem_nfee_comm_1:avs_0_rmap_write_i
	wire   [31:0] mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_writedata;                      // mm_interconnect_1:rmap_mem_nfee_comm_1_avalon_rmap_slave_0_writedata -> rmap_mem_nfee_comm_1:avs_0_rmap_writedata_i
	wire   [31:0] mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_readdata;                       // rmap_mem_nfee_comm_2:avs_0_rmap_readdata_o -> mm_interconnect_1:rmap_mem_nfee_comm_2_avalon_rmap_slave_0_readdata
	wire          mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_waitrequest;                    // rmap_mem_nfee_comm_2:avs_0_rmap_waitrequest_o -> mm_interconnect_1:rmap_mem_nfee_comm_2_avalon_rmap_slave_0_waitrequest
	wire   [11:0] mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_address;                        // mm_interconnect_1:rmap_mem_nfee_comm_2_avalon_rmap_slave_0_address -> rmap_mem_nfee_comm_2:avs_0_rmap_address_i
	wire          mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_read;                           // mm_interconnect_1:rmap_mem_nfee_comm_2_avalon_rmap_slave_0_read -> rmap_mem_nfee_comm_2:avs_0_rmap_read_i
	wire    [3:0] mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_byteenable;                     // mm_interconnect_1:rmap_mem_nfee_comm_2_avalon_rmap_slave_0_byteenable -> rmap_mem_nfee_comm_2:avs_0_rmap_byteenable_i
	wire          mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_write;                          // mm_interconnect_1:rmap_mem_nfee_comm_2_avalon_rmap_slave_0_write -> rmap_mem_nfee_comm_2:avs_0_rmap_write_i
	wire   [31:0] mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_writedata;                      // mm_interconnect_1:rmap_mem_nfee_comm_2_avalon_rmap_slave_0_writedata -> rmap_mem_nfee_comm_2:avs_0_rmap_writedata_i
	wire   [31:0] mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_readdata;                       // rmap_mem_nfee_comm_3:avs_0_rmap_readdata_o -> mm_interconnect_1:rmap_mem_nfee_comm_3_avalon_rmap_slave_0_readdata
	wire          mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_waitrequest;                    // rmap_mem_nfee_comm_3:avs_0_rmap_waitrequest_o -> mm_interconnect_1:rmap_mem_nfee_comm_3_avalon_rmap_slave_0_waitrequest
	wire   [11:0] mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_address;                        // mm_interconnect_1:rmap_mem_nfee_comm_3_avalon_rmap_slave_0_address -> rmap_mem_nfee_comm_3:avs_0_rmap_address_i
	wire          mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_read;                           // mm_interconnect_1:rmap_mem_nfee_comm_3_avalon_rmap_slave_0_read -> rmap_mem_nfee_comm_3:avs_0_rmap_read_i
	wire    [3:0] mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_byteenable;                     // mm_interconnect_1:rmap_mem_nfee_comm_3_avalon_rmap_slave_0_byteenable -> rmap_mem_nfee_comm_3:avs_0_rmap_byteenable_i
	wire          mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_write;                          // mm_interconnect_1:rmap_mem_nfee_comm_3_avalon_rmap_slave_0_write -> rmap_mem_nfee_comm_3:avs_0_rmap_write_i
	wire   [31:0] mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_writedata;                      // mm_interconnect_1:rmap_mem_nfee_comm_3_avalon_rmap_slave_0_writedata -> rmap_mem_nfee_comm_3:avs_0_rmap_writedata_i
	wire   [31:0] mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_readdata;                       // rmap_mem_nfee_comm_4:avs_0_rmap_readdata_o -> mm_interconnect_1:rmap_mem_nfee_comm_4_avalon_rmap_slave_0_readdata
	wire          mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_waitrequest;                    // rmap_mem_nfee_comm_4:avs_0_rmap_waitrequest_o -> mm_interconnect_1:rmap_mem_nfee_comm_4_avalon_rmap_slave_0_waitrequest
	wire   [11:0] mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_address;                        // mm_interconnect_1:rmap_mem_nfee_comm_4_avalon_rmap_slave_0_address -> rmap_mem_nfee_comm_4:avs_0_rmap_address_i
	wire          mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_read;                           // mm_interconnect_1:rmap_mem_nfee_comm_4_avalon_rmap_slave_0_read -> rmap_mem_nfee_comm_4:avs_0_rmap_read_i
	wire    [3:0] mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_byteenable;                     // mm_interconnect_1:rmap_mem_nfee_comm_4_avalon_rmap_slave_0_byteenable -> rmap_mem_nfee_comm_4:avs_0_rmap_byteenable_i
	wire          mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_write;                          // mm_interconnect_1:rmap_mem_nfee_comm_4_avalon_rmap_slave_0_write -> rmap_mem_nfee_comm_4:avs_0_rmap_write_i
	wire   [31:0] mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_writedata;                      // mm_interconnect_1:rmap_mem_nfee_comm_4_avalon_rmap_slave_0_writedata -> rmap_mem_nfee_comm_4:avs_0_rmap_writedata_i
	wire   [31:0] mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_readdata;                       // rmap_mem_nfee_comm_5:avs_0_rmap_readdata_o -> mm_interconnect_1:rmap_mem_nfee_comm_5_avalon_rmap_slave_0_readdata
	wire          mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_waitrequest;                    // rmap_mem_nfee_comm_5:avs_0_rmap_waitrequest_o -> mm_interconnect_1:rmap_mem_nfee_comm_5_avalon_rmap_slave_0_waitrequest
	wire   [11:0] mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_address;                        // mm_interconnect_1:rmap_mem_nfee_comm_5_avalon_rmap_slave_0_address -> rmap_mem_nfee_comm_5:avs_0_rmap_address_i
	wire          mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_read;                           // mm_interconnect_1:rmap_mem_nfee_comm_5_avalon_rmap_slave_0_read -> rmap_mem_nfee_comm_5:avs_0_rmap_read_i
	wire    [3:0] mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_byteenable;                     // mm_interconnect_1:rmap_mem_nfee_comm_5_avalon_rmap_slave_0_byteenable -> rmap_mem_nfee_comm_5:avs_0_rmap_byteenable_i
	wire          mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_write;                          // mm_interconnect_1:rmap_mem_nfee_comm_5_avalon_rmap_slave_0_write -> rmap_mem_nfee_comm_5:avs_0_rmap_write_i
	wire   [31:0] mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_writedata;                      // mm_interconnect_1:rmap_mem_nfee_comm_5_avalon_rmap_slave_0_writedata -> rmap_mem_nfee_comm_5:avs_0_rmap_writedata_i
	wire   [31:0] mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_readdata;                       // rmap_mem_nfee_comm_6:avs_0_rmap_readdata_o -> mm_interconnect_1:rmap_mem_nfee_comm_6_avalon_rmap_slave_0_readdata
	wire          mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_waitrequest;                    // rmap_mem_nfee_comm_6:avs_0_rmap_waitrequest_o -> mm_interconnect_1:rmap_mem_nfee_comm_6_avalon_rmap_slave_0_waitrequest
	wire   [11:0] mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_address;                        // mm_interconnect_1:rmap_mem_nfee_comm_6_avalon_rmap_slave_0_address -> rmap_mem_nfee_comm_6:avs_0_rmap_address_i
	wire          mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_read;                           // mm_interconnect_1:rmap_mem_nfee_comm_6_avalon_rmap_slave_0_read -> rmap_mem_nfee_comm_6:avs_0_rmap_read_i
	wire    [3:0] mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_byteenable;                     // mm_interconnect_1:rmap_mem_nfee_comm_6_avalon_rmap_slave_0_byteenable -> rmap_mem_nfee_comm_6:avs_0_rmap_byteenable_i
	wire          mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_write;                          // mm_interconnect_1:rmap_mem_nfee_comm_6_avalon_rmap_slave_0_write -> rmap_mem_nfee_comm_6:avs_0_rmap_write_i
	wire   [31:0] mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_writedata;                      // mm_interconnect_1:rmap_mem_nfee_comm_6_avalon_rmap_slave_0_writedata -> rmap_mem_nfee_comm_6:avs_0_rmap_writedata_i
	wire   [31:0] mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_readdata;                                // FTDI_USB3_0:avalon_slave_config_readdata -> mm_interconnect_1:FTDI_USB3_0_avalon_slave_config_readdata
	wire          mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_waitrequest;                             // FTDI_USB3_0:avalon_slave_config_waitrequest -> mm_interconnect_1:FTDI_USB3_0_avalon_slave_config_waitrequest
	wire    [7:0] mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_address;                                 // mm_interconnect_1:FTDI_USB3_0_avalon_slave_config_address -> FTDI_USB3_0:avalon_slave_config_address
	wire          mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_read;                                    // mm_interconnect_1:FTDI_USB3_0_avalon_slave_config_read -> FTDI_USB3_0:avalon_slave_config_read
	wire    [3:0] mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_byteenable;                              // mm_interconnect_1:FTDI_USB3_0_avalon_slave_config_byteenable -> FTDI_USB3_0:avalon_slave_config_byteenable
	wire          mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_write;                                   // mm_interconnect_1:FTDI_USB3_0_avalon_slave_config_write -> FTDI_USB3_0:avalon_slave_config_write
	wire   [31:0] mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_writedata;                               // mm_interconnect_1:FTDI_USB3_0_avalon_slave_config_writedata -> FTDI_USB3_0:avalon_slave_config_writedata
	wire   [31:0] mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_readdata;                   // COMM_Pedreiro_v1_01_1:avalon_slave_windowing_readdata -> mm_interconnect_1:COMM_Pedreiro_v1_01_1_avalon_slave_windowing_readdata
	wire          mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_waitrequest;                // COMM_Pedreiro_v1_01_1:avalon_slave_windowing_waitrequest -> mm_interconnect_1:COMM_Pedreiro_v1_01_1_avalon_slave_windowing_waitrequest
	wire    [7:0] mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_address;                    // mm_interconnect_1:COMM_Pedreiro_v1_01_1_avalon_slave_windowing_address -> COMM_Pedreiro_v1_01_1:avalon_slave_windowing_address
	wire          mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_read;                       // mm_interconnect_1:COMM_Pedreiro_v1_01_1_avalon_slave_windowing_read -> COMM_Pedreiro_v1_01_1:avalon_slave_windowing_read
	wire    [3:0] mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_byteenable;                 // mm_interconnect_1:COMM_Pedreiro_v1_01_1_avalon_slave_windowing_byteenable -> COMM_Pedreiro_v1_01_1:avalon_slave_windowing_byteenable
	wire          mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_write;                      // mm_interconnect_1:COMM_Pedreiro_v1_01_1_avalon_slave_windowing_write -> COMM_Pedreiro_v1_01_1:avalon_slave_windowing_write
	wire   [31:0] mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_writedata;                  // mm_interconnect_1:COMM_Pedreiro_v1_01_1_avalon_slave_windowing_writedata -> COMM_Pedreiro_v1_01_1:avalon_slave_windowing_writedata
	wire   [31:0] mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_readdata;                   // COMM_Pedreiro_v1_01_2:avalon_slave_windowing_readdata -> mm_interconnect_1:COMM_Pedreiro_v1_01_2_avalon_slave_windowing_readdata
	wire          mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_waitrequest;                // COMM_Pedreiro_v1_01_2:avalon_slave_windowing_waitrequest -> mm_interconnect_1:COMM_Pedreiro_v1_01_2_avalon_slave_windowing_waitrequest
	wire    [7:0] mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_address;                    // mm_interconnect_1:COMM_Pedreiro_v1_01_2_avalon_slave_windowing_address -> COMM_Pedreiro_v1_01_2:avalon_slave_windowing_address
	wire          mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_read;                       // mm_interconnect_1:COMM_Pedreiro_v1_01_2_avalon_slave_windowing_read -> COMM_Pedreiro_v1_01_2:avalon_slave_windowing_read
	wire    [3:0] mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_byteenable;                 // mm_interconnect_1:COMM_Pedreiro_v1_01_2_avalon_slave_windowing_byteenable -> COMM_Pedreiro_v1_01_2:avalon_slave_windowing_byteenable
	wire          mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_write;                      // mm_interconnect_1:COMM_Pedreiro_v1_01_2_avalon_slave_windowing_write -> COMM_Pedreiro_v1_01_2:avalon_slave_windowing_write
	wire   [31:0] mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_writedata;                  // mm_interconnect_1:COMM_Pedreiro_v1_01_2_avalon_slave_windowing_writedata -> COMM_Pedreiro_v1_01_2:avalon_slave_windowing_writedata
	wire   [31:0] mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_readdata;                   // COMM_Pedreiro_v1_01_3:avalon_slave_windowing_readdata -> mm_interconnect_1:COMM_Pedreiro_v1_01_3_avalon_slave_windowing_readdata
	wire          mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_waitrequest;                // COMM_Pedreiro_v1_01_3:avalon_slave_windowing_waitrequest -> mm_interconnect_1:COMM_Pedreiro_v1_01_3_avalon_slave_windowing_waitrequest
	wire    [7:0] mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_address;                    // mm_interconnect_1:COMM_Pedreiro_v1_01_3_avalon_slave_windowing_address -> COMM_Pedreiro_v1_01_3:avalon_slave_windowing_address
	wire          mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_read;                       // mm_interconnect_1:COMM_Pedreiro_v1_01_3_avalon_slave_windowing_read -> COMM_Pedreiro_v1_01_3:avalon_slave_windowing_read
	wire    [3:0] mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_byteenable;                 // mm_interconnect_1:COMM_Pedreiro_v1_01_3_avalon_slave_windowing_byteenable -> COMM_Pedreiro_v1_01_3:avalon_slave_windowing_byteenable
	wire          mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_write;                      // mm_interconnect_1:COMM_Pedreiro_v1_01_3_avalon_slave_windowing_write -> COMM_Pedreiro_v1_01_3:avalon_slave_windowing_write
	wire   [31:0] mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_writedata;                  // mm_interconnect_1:COMM_Pedreiro_v1_01_3_avalon_slave_windowing_writedata -> COMM_Pedreiro_v1_01_3:avalon_slave_windowing_writedata
	wire   [31:0] mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_readdata;                   // COMM_Pedreiro_v1_01_4:avalon_slave_windowing_readdata -> mm_interconnect_1:COMM_Pedreiro_v1_01_4_avalon_slave_windowing_readdata
	wire          mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_waitrequest;                // COMM_Pedreiro_v1_01_4:avalon_slave_windowing_waitrequest -> mm_interconnect_1:COMM_Pedreiro_v1_01_4_avalon_slave_windowing_waitrequest
	wire    [7:0] mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_address;                    // mm_interconnect_1:COMM_Pedreiro_v1_01_4_avalon_slave_windowing_address -> COMM_Pedreiro_v1_01_4:avalon_slave_windowing_address
	wire          mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_read;                       // mm_interconnect_1:COMM_Pedreiro_v1_01_4_avalon_slave_windowing_read -> COMM_Pedreiro_v1_01_4:avalon_slave_windowing_read
	wire    [3:0] mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_byteenable;                 // mm_interconnect_1:COMM_Pedreiro_v1_01_4_avalon_slave_windowing_byteenable -> COMM_Pedreiro_v1_01_4:avalon_slave_windowing_byteenable
	wire          mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_write;                      // mm_interconnect_1:COMM_Pedreiro_v1_01_4_avalon_slave_windowing_write -> COMM_Pedreiro_v1_01_4:avalon_slave_windowing_write
	wire   [31:0] mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_writedata;                  // mm_interconnect_1:COMM_Pedreiro_v1_01_4_avalon_slave_windowing_writedata -> COMM_Pedreiro_v1_01_4:avalon_slave_windowing_writedata
	wire   [31:0] mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_readdata;                   // COMM_Pedreiro_v1_01_5:avalon_slave_windowing_readdata -> mm_interconnect_1:COMM_Pedreiro_v1_01_5_avalon_slave_windowing_readdata
	wire          mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_waitrequest;                // COMM_Pedreiro_v1_01_5:avalon_slave_windowing_waitrequest -> mm_interconnect_1:COMM_Pedreiro_v1_01_5_avalon_slave_windowing_waitrequest
	wire    [7:0] mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_address;                    // mm_interconnect_1:COMM_Pedreiro_v1_01_5_avalon_slave_windowing_address -> COMM_Pedreiro_v1_01_5:avalon_slave_windowing_address
	wire          mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_read;                       // mm_interconnect_1:COMM_Pedreiro_v1_01_5_avalon_slave_windowing_read -> COMM_Pedreiro_v1_01_5:avalon_slave_windowing_read
	wire    [3:0] mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_byteenable;                 // mm_interconnect_1:COMM_Pedreiro_v1_01_5_avalon_slave_windowing_byteenable -> COMM_Pedreiro_v1_01_5:avalon_slave_windowing_byteenable
	wire          mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_write;                      // mm_interconnect_1:COMM_Pedreiro_v1_01_5_avalon_slave_windowing_write -> COMM_Pedreiro_v1_01_5:avalon_slave_windowing_write
	wire   [31:0] mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_writedata;                  // mm_interconnect_1:COMM_Pedreiro_v1_01_5_avalon_slave_windowing_writedata -> COMM_Pedreiro_v1_01_5:avalon_slave_windowing_writedata
	wire   [31:0] mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_readdata;                   // COMM_Pedreiro_v1_01_6:avalon_slave_windowing_readdata -> mm_interconnect_1:COMM_Pedreiro_v1_01_6_avalon_slave_windowing_readdata
	wire          mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_waitrequest;                // COMM_Pedreiro_v1_01_6:avalon_slave_windowing_waitrequest -> mm_interconnect_1:COMM_Pedreiro_v1_01_6_avalon_slave_windowing_waitrequest
	wire    [7:0] mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_address;                    // mm_interconnect_1:COMM_Pedreiro_v1_01_6_avalon_slave_windowing_address -> COMM_Pedreiro_v1_01_6:avalon_slave_windowing_address
	wire          mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_read;                       // mm_interconnect_1:COMM_Pedreiro_v1_01_6_avalon_slave_windowing_read -> COMM_Pedreiro_v1_01_6:avalon_slave_windowing_read
	wire    [3:0] mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_byteenable;                 // mm_interconnect_1:COMM_Pedreiro_v1_01_6_avalon_slave_windowing_byteenable -> COMM_Pedreiro_v1_01_6:avalon_slave_windowing_byteenable
	wire          mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_write;                      // mm_interconnect_1:COMM_Pedreiro_v1_01_6_avalon_slave_windowing_write -> COMM_Pedreiro_v1_01_6:avalon_slave_windowing_write
	wire   [31:0] mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_writedata;                  // mm_interconnect_1:COMM_Pedreiro_v1_01_6_avalon_slave_windowing_writedata -> COMM_Pedreiro_v1_01_6:avalon_slave_windowing_writedata
	wire   [63:0] mm_interconnect_1_ddr2_address_span_extender_cntl_readdata;                                // ddr2_address_span_extender:avs_cntl_readdata -> mm_interconnect_1:ddr2_address_span_extender_cntl_readdata
	wire          mm_interconnect_1_ddr2_address_span_extender_cntl_read;                                    // mm_interconnect_1:ddr2_address_span_extender_cntl_read -> ddr2_address_span_extender:avs_cntl_read
	wire    [7:0] mm_interconnect_1_ddr2_address_span_extender_cntl_byteenable;                              // mm_interconnect_1:ddr2_address_span_extender_cntl_byteenable -> ddr2_address_span_extender:avs_cntl_byteenable
	wire          mm_interconnect_1_ddr2_address_span_extender_cntl_write;                                   // mm_interconnect_1:ddr2_address_span_extender_cntl_write -> ddr2_address_span_extender:avs_cntl_write
	wire   [63:0] mm_interconnect_1_ddr2_address_span_extender_cntl_writedata;                               // mm_interconnect_1:ddr2_address_span_extender_cntl_writedata -> ddr2_address_span_extender:avs_cntl_writedata
	wire   [31:0] mm_interconnect_1_sysid_qsys_control_slave_readdata;                                       // sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	wire    [0:0] mm_interconnect_1_sysid_qsys_control_slave_address;                                        // mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire   [31:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata;                                   // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_readdata
	wire          mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest;                                // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_waitrequest
	wire          mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess;                                // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address;                                    // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire          mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read;                                       // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire    [3:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable;                                 // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire          mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write;                                      // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire   [31:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata;                                  // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire   [31:0] mm_interconnect_1_clock_bridge_afi_50_s0_readdata;                                         // clock_bridge_afi_50:s0_readdata -> mm_interconnect_1:clock_bridge_afi_50_s0_readdata
	wire          mm_interconnect_1_clock_bridge_afi_50_s0_waitrequest;                                      // clock_bridge_afi_50:s0_waitrequest -> mm_interconnect_1:clock_bridge_afi_50_s0_waitrequest
	wire          mm_interconnect_1_clock_bridge_afi_50_s0_debugaccess;                                      // mm_interconnect_1:clock_bridge_afi_50_s0_debugaccess -> clock_bridge_afi_50:s0_debugaccess
	wire   [11:0] mm_interconnect_1_clock_bridge_afi_50_s0_address;                                          // mm_interconnect_1:clock_bridge_afi_50_s0_address -> clock_bridge_afi_50:s0_address
	wire          mm_interconnect_1_clock_bridge_afi_50_s0_read;                                             // mm_interconnect_1:clock_bridge_afi_50_s0_read -> clock_bridge_afi_50:s0_read
	wire    [3:0] mm_interconnect_1_clock_bridge_afi_50_s0_byteenable;                                       // mm_interconnect_1:clock_bridge_afi_50_s0_byteenable -> clock_bridge_afi_50:s0_byteenable
	wire          mm_interconnect_1_clock_bridge_afi_50_s0_readdatavalid;                                    // clock_bridge_afi_50:s0_readdatavalid -> mm_interconnect_1:clock_bridge_afi_50_s0_readdatavalid
	wire          mm_interconnect_1_clock_bridge_afi_50_s0_write;                                            // mm_interconnect_1:clock_bridge_afi_50_s0_write -> clock_bridge_afi_50:s0_write
	wire   [31:0] mm_interconnect_1_clock_bridge_afi_50_s0_writedata;                                        // mm_interconnect_1:clock_bridge_afi_50_s0_writedata -> clock_bridge_afi_50:s0_writedata
	wire    [0:0] mm_interconnect_1_clock_bridge_afi_50_s0_burstcount;                                       // mm_interconnect_1:clock_bridge_afi_50_s0_burstcount -> clock_bridge_afi_50:s0_burstcount
	wire          mm_interconnect_1_onchip_memory_s1_chipselect;                                             // mm_interconnect_1:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire   [31:0] mm_interconnect_1_onchip_memory_s1_readdata;                                               // onchip_memory:readdata -> mm_interconnect_1:onchip_memory_s1_readdata
	wire   [17:0] mm_interconnect_1_onchip_memory_s1_address;                                                // mm_interconnect_1:onchip_memory_s1_address -> onchip_memory:address
	wire    [3:0] mm_interconnect_1_onchip_memory_s1_byteenable;                                             // mm_interconnect_1:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire          mm_interconnect_1_onchip_memory_s1_write;                                                  // mm_interconnect_1:onchip_memory_s1_write -> onchip_memory:write
	wire   [31:0] mm_interconnect_1_onchip_memory_s1_writedata;                                              // mm_interconnect_1:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire          mm_interconnect_1_onchip_memory_s1_clken;                                                  // mm_interconnect_1:onchip_memory_s1_clken -> onchip_memory:clken
	wire   [15:0] mm_interconnect_1_ext_flash_uas_readdata;                                                  // ext_flash:uas_readdata -> mm_interconnect_1:ext_flash_uas_readdata
	wire          mm_interconnect_1_ext_flash_uas_waitrequest;                                               // ext_flash:uas_waitrequest -> mm_interconnect_1:ext_flash_uas_waitrequest
	wire          mm_interconnect_1_ext_flash_uas_debugaccess;                                               // mm_interconnect_1:ext_flash_uas_debugaccess -> ext_flash:uas_debugaccess
	wire   [25:0] mm_interconnect_1_ext_flash_uas_address;                                                   // mm_interconnect_1:ext_flash_uas_address -> ext_flash:uas_address
	wire          mm_interconnect_1_ext_flash_uas_read;                                                      // mm_interconnect_1:ext_flash_uas_read -> ext_flash:uas_read
	wire    [1:0] mm_interconnect_1_ext_flash_uas_byteenable;                                                // mm_interconnect_1:ext_flash_uas_byteenable -> ext_flash:uas_byteenable
	wire          mm_interconnect_1_ext_flash_uas_readdatavalid;                                             // ext_flash:uas_readdatavalid -> mm_interconnect_1:ext_flash_uas_readdatavalid
	wire          mm_interconnect_1_ext_flash_uas_lock;                                                      // mm_interconnect_1:ext_flash_uas_lock -> ext_flash:uas_lock
	wire          mm_interconnect_1_ext_flash_uas_write;                                                     // mm_interconnect_1:ext_flash_uas_write -> ext_flash:uas_write
	wire   [15:0] mm_interconnect_1_ext_flash_uas_writedata;                                                 // mm_interconnect_1:ext_flash_uas_writedata -> ext_flash:uas_writedata
	wire    [1:0] mm_interconnect_1_ext_flash_uas_burstcount;                                                // mm_interconnect_1:ext_flash_uas_burstcount -> ext_flash:uas_burstcount
	wire   [31:0] mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdata;                      // ddr2_address_span_extender:avs_s0_readdata -> mm_interconnect_1:ddr2_address_span_extender_windowed_slave_readdata
	wire          mm_interconnect_1_ddr2_address_span_extender_windowed_slave_waitrequest;                   // ddr2_address_span_extender:avs_s0_waitrequest -> mm_interconnect_1:ddr2_address_span_extender_windowed_slave_waitrequest
	wire   [28:0] mm_interconnect_1_ddr2_address_span_extender_windowed_slave_address;                       // mm_interconnect_1:ddr2_address_span_extender_windowed_slave_address -> ddr2_address_span_extender:avs_s0_address
	wire          mm_interconnect_1_ddr2_address_span_extender_windowed_slave_read;                          // mm_interconnect_1:ddr2_address_span_extender_windowed_slave_read -> ddr2_address_span_extender:avs_s0_read
	wire    [3:0] mm_interconnect_1_ddr2_address_span_extender_windowed_slave_byteenable;                    // mm_interconnect_1:ddr2_address_span_extender_windowed_slave_byteenable -> ddr2_address_span_extender:avs_s0_byteenable
	wire          mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdatavalid;                 // ddr2_address_span_extender:avs_s0_readdatavalid -> mm_interconnect_1:ddr2_address_span_extender_windowed_slave_readdatavalid
	wire          mm_interconnect_1_ddr2_address_span_extender_windowed_slave_write;                         // mm_interconnect_1:ddr2_address_span_extender_windowed_slave_write -> ddr2_address_span_extender:avs_s0_write
	wire   [31:0] mm_interconnect_1_ddr2_address_span_extender_windowed_slave_writedata;                     // mm_interconnect_1:ddr2_address_span_extender_windowed_slave_writedata -> ddr2_address_span_extender:avs_s0_writedata
	wire    [7:0] mm_interconnect_1_ddr2_address_span_extender_windowed_slave_burstcount;                    // mm_interconnect_1:ddr2_address_span_extender_windowed_slave_burstcount -> ddr2_address_span_extender:avs_s0_burstcount
	wire          clock_bridge_afi_50_m0_waitrequest;                                                        // mm_interconnect_2:clock_bridge_afi_50_m0_waitrequest -> clock_bridge_afi_50:m0_waitrequest
	wire   [31:0] clock_bridge_afi_50_m0_readdata;                                                           // mm_interconnect_2:clock_bridge_afi_50_m0_readdata -> clock_bridge_afi_50:m0_readdata
	wire          clock_bridge_afi_50_m0_debugaccess;                                                        // clock_bridge_afi_50:m0_debugaccess -> mm_interconnect_2:clock_bridge_afi_50_m0_debugaccess
	wire   [11:0] clock_bridge_afi_50_m0_address;                                                            // clock_bridge_afi_50:m0_address -> mm_interconnect_2:clock_bridge_afi_50_m0_address
	wire          clock_bridge_afi_50_m0_read;                                                               // clock_bridge_afi_50:m0_read -> mm_interconnect_2:clock_bridge_afi_50_m0_read
	wire    [3:0] clock_bridge_afi_50_m0_byteenable;                                                         // clock_bridge_afi_50:m0_byteenable -> mm_interconnect_2:clock_bridge_afi_50_m0_byteenable
	wire          clock_bridge_afi_50_m0_readdatavalid;                                                      // mm_interconnect_2:clock_bridge_afi_50_m0_readdatavalid -> clock_bridge_afi_50:m0_readdatavalid
	wire   [31:0] clock_bridge_afi_50_m0_writedata;                                                          // clock_bridge_afi_50:m0_writedata -> mm_interconnect_2:clock_bridge_afi_50_m0_writedata
	wire          clock_bridge_afi_50_m0_write;                                                              // clock_bridge_afi_50:m0_write -> mm_interconnect_2:clock_bridge_afi_50_m0_write
	wire    [0:0] clock_bridge_afi_50_m0_burstcount;                                                         // clock_bridge_afi_50:m0_burstcount -> mm_interconnect_2:clock_bridge_afi_50_m0_burstcount
	wire   [31:0] mm_interconnect_2_sync_avalon_mm_slave_readdata;                                           // sync:avalon_slave_readdata_o -> mm_interconnect_2:sync_avalon_mm_slave_readdata
	wire          mm_interconnect_2_sync_avalon_mm_slave_waitrequest;                                        // sync:avalon_slave_waitrequest_o -> mm_interconnect_2:sync_avalon_mm_slave_waitrequest
	wire    [7:0] mm_interconnect_2_sync_avalon_mm_slave_address;                                            // mm_interconnect_2:sync_avalon_mm_slave_address -> sync:avalon_slave_address_i
	wire          mm_interconnect_2_sync_avalon_mm_slave_read;                                               // mm_interconnect_2:sync_avalon_mm_slave_read -> sync:avalon_slave_read_i
	wire    [3:0] mm_interconnect_2_sync_avalon_mm_slave_byteenable;                                         // mm_interconnect_2:sync_avalon_mm_slave_byteenable -> sync:avalon_slave_byteenable_i
	wire          mm_interconnect_2_sync_avalon_mm_slave_write;                                              // mm_interconnect_2:sync_avalon_mm_slave_write -> sync:avalon_slave_write_i
	wire   [31:0] mm_interconnect_2_sync_avalon_mm_slave_writedata;                                          // mm_interconnect_2:sync_avalon_mm_slave_writedata -> sync:avalon_slave_writedata_i
	wire   [31:0] mm_interconnect_2_rst_controller_avalon_rst_controller_slave_readdata;                     // rst_controller:avalon_slave_rst_controller_readdata -> mm_interconnect_2:rst_controller_avalon_rst_controller_slave_readdata
	wire          mm_interconnect_2_rst_controller_avalon_rst_controller_slave_waitrequest;                  // rst_controller:avalon_slave_rst_controller_waitrequest -> mm_interconnect_2:rst_controller_avalon_rst_controller_slave_waitrequest
	wire    [3:0] mm_interconnect_2_rst_controller_avalon_rst_controller_slave_address;                      // mm_interconnect_2:rst_controller_avalon_rst_controller_slave_address -> rst_controller:avalon_slave_rst_controller_address
	wire          mm_interconnect_2_rst_controller_avalon_rst_controller_slave_read;                         // mm_interconnect_2:rst_controller_avalon_rst_controller_slave_read -> rst_controller:avalon_slave_rst_controller_read
	wire          mm_interconnect_2_rst_controller_avalon_rst_controller_slave_write;                        // mm_interconnect_2:rst_controller_avalon_rst_controller_slave_write -> rst_controller:avalon_slave_rst_controller_write
	wire   [31:0] mm_interconnect_2_rst_controller_avalon_rst_controller_slave_writedata;                    // mm_interconnect_2:rst_controller_avalon_rst_controller_slave_writedata -> rst_controller:avalon_slave_rst_controller_writedata
	wire          mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect;     // mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_chip_select
	wire   [31:0] mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata;       // Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_readdata -> mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata
	wire          mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest;    // Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_waitrequest -> mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest
	wire    [7:0] mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address;        // mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_address
	wire          mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read;           // mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_read
	wire    [3:0] mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable;     // mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_byteenable
	wire          mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write;          // mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_write
	wire   [31:0] mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata;      // mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_writedata
	wire          mm_interconnect_2_m1_ddr2_i2c_sda_s1_chipselect;                                           // mm_interconnect_2:m1_ddr2_i2c_sda_s1_chipselect -> m1_ddr2_i2c_sda:chipselect
	wire   [31:0] mm_interconnect_2_m1_ddr2_i2c_sda_s1_readdata;                                             // m1_ddr2_i2c_sda:readdata -> mm_interconnect_2:m1_ddr2_i2c_sda_s1_readdata
	wire    [1:0] mm_interconnect_2_m1_ddr2_i2c_sda_s1_address;                                              // mm_interconnect_2:m1_ddr2_i2c_sda_s1_address -> m1_ddr2_i2c_sda:address
	wire          mm_interconnect_2_m1_ddr2_i2c_sda_s1_write;                                                // mm_interconnect_2:m1_ddr2_i2c_sda_s1_write -> m1_ddr2_i2c_sda:write_n
	wire   [31:0] mm_interconnect_2_m1_ddr2_i2c_sda_s1_writedata;                                            // mm_interconnect_2:m1_ddr2_i2c_sda_s1_writedata -> m1_ddr2_i2c_sda:writedata
	wire          mm_interconnect_2_m1_ddr2_i2c_scl_s1_chipselect;                                           // mm_interconnect_2:m1_ddr2_i2c_scl_s1_chipselect -> m1_ddr2_i2c_scl:chipselect
	wire   [31:0] mm_interconnect_2_m1_ddr2_i2c_scl_s1_readdata;                                             // m1_ddr2_i2c_scl:readdata -> mm_interconnect_2:m1_ddr2_i2c_scl_s1_readdata
	wire    [1:0] mm_interconnect_2_m1_ddr2_i2c_scl_s1_address;                                              // mm_interconnect_2:m1_ddr2_i2c_scl_s1_address -> m1_ddr2_i2c_scl:address
	wire          mm_interconnect_2_m1_ddr2_i2c_scl_s1_write;                                                // mm_interconnect_2:m1_ddr2_i2c_scl_s1_write -> m1_ddr2_i2c_scl:write_n
	wire   [31:0] mm_interconnect_2_m1_ddr2_i2c_scl_s1_writedata;                                            // mm_interconnect_2:m1_ddr2_i2c_scl_s1_writedata -> m1_ddr2_i2c_scl:writedata
	wire   [31:0] mm_interconnect_2_pio_button_s1_readdata;                                                  // pio_BUTTON:readdata -> mm_interconnect_2:pio_BUTTON_s1_readdata
	wire    [1:0] mm_interconnect_2_pio_button_s1_address;                                                   // mm_interconnect_2:pio_BUTTON_s1_address -> pio_BUTTON:address
	wire          mm_interconnect_2_pio_led_s1_chipselect;                                                   // mm_interconnect_2:pio_LED_s1_chipselect -> pio_LED:chipselect
	wire   [31:0] mm_interconnect_2_pio_led_s1_readdata;                                                     // pio_LED:readdata -> mm_interconnect_2:pio_LED_s1_readdata
	wire    [1:0] mm_interconnect_2_pio_led_s1_address;                                                      // mm_interconnect_2:pio_LED_s1_address -> pio_LED:address
	wire          mm_interconnect_2_pio_led_s1_write;                                                        // mm_interconnect_2:pio_LED_s1_write -> pio_LED:write_n
	wire   [31:0] mm_interconnect_2_pio_led_s1_writedata;                                                    // mm_interconnect_2:pio_LED_s1_writedata -> pio_LED:writedata
	wire          mm_interconnect_2_timer_1ms_s1_chipselect;                                                 // mm_interconnect_2:timer_1ms_s1_chipselect -> timer_1ms:chipselect
	wire   [15:0] mm_interconnect_2_timer_1ms_s1_readdata;                                                   // timer_1ms:readdata -> mm_interconnect_2:timer_1ms_s1_readdata
	wire    [2:0] mm_interconnect_2_timer_1ms_s1_address;                                                    // mm_interconnect_2:timer_1ms_s1_address -> timer_1ms:address
	wire          mm_interconnect_2_timer_1ms_s1_write;                                                      // mm_interconnect_2:timer_1ms_s1_write -> timer_1ms:write_n
	wire   [15:0] mm_interconnect_2_timer_1ms_s1_writedata;                                                  // mm_interconnect_2:timer_1ms_s1_writedata -> timer_1ms:writedata
	wire   [31:0] mm_interconnect_2_pio_dip_s1_readdata;                                                     // pio_DIP:readdata -> mm_interconnect_2:pio_DIP_s1_readdata
	wire    [1:0] mm_interconnect_2_pio_dip_s1_address;                                                      // mm_interconnect_2:pio_DIP_s1_address -> pio_DIP:address
	wire          mm_interconnect_2_timer_1us_s1_chipselect;                                                 // mm_interconnect_2:timer_1us_s1_chipselect -> timer_1us:chipselect
	wire   [15:0] mm_interconnect_2_timer_1us_s1_readdata;                                                   // timer_1us:readdata -> mm_interconnect_2:timer_1us_s1_readdata
	wire    [2:0] mm_interconnect_2_timer_1us_s1_address;                                                    // mm_interconnect_2:timer_1us_s1_address -> timer_1us:address
	wire          mm_interconnect_2_timer_1us_s1_write;                                                      // mm_interconnect_2:timer_1us_s1_write -> timer_1us:write_n
	wire   [15:0] mm_interconnect_2_timer_1us_s1_writedata;                                                  // mm_interconnect_2:timer_1us_s1_writedata -> timer_1us:writedata
	wire   [31:0] mm_interconnect_2_pio_ext_s1_readdata;                                                     // pio_EXT:readdata -> mm_interconnect_2:pio_EXT_s1_readdata
	wire    [1:0] mm_interconnect_2_pio_ext_s1_address;                                                      // mm_interconnect_2:pio_EXT_s1_address -> pio_EXT:address
	wire   [31:0] mm_interconnect_2_sd_card_wp_n_s1_readdata;                                                // sd_card_wp_n:readdata -> mm_interconnect_2:sd_card_wp_n_s1_readdata
	wire    [1:0] mm_interconnect_2_sd_card_wp_n_s1_address;                                                 // mm_interconnect_2:sd_card_wp_n_s1_address -> sd_card_wp_n:address
	wire          mm_interconnect_2_temp_scl_s1_chipselect;                                                  // mm_interconnect_2:temp_scl_s1_chipselect -> temp_scl:chipselect
	wire   [31:0] mm_interconnect_2_temp_scl_s1_readdata;                                                    // temp_scl:readdata -> mm_interconnect_2:temp_scl_s1_readdata
	wire    [1:0] mm_interconnect_2_temp_scl_s1_address;                                                     // mm_interconnect_2:temp_scl_s1_address -> temp_scl:address
	wire          mm_interconnect_2_temp_scl_s1_write;                                                       // mm_interconnect_2:temp_scl_s1_write -> temp_scl:write_n
	wire   [31:0] mm_interconnect_2_temp_scl_s1_writedata;                                                   // mm_interconnect_2:temp_scl_s1_writedata -> temp_scl:writedata
	wire          mm_interconnect_2_temp_sda_s1_chipselect;                                                  // mm_interconnect_2:temp_sda_s1_chipselect -> temp_sda:chipselect
	wire   [31:0] mm_interconnect_2_temp_sda_s1_readdata;                                                    // temp_sda:readdata -> mm_interconnect_2:temp_sda_s1_readdata
	wire    [1:0] mm_interconnect_2_temp_sda_s1_address;                                                     // mm_interconnect_2:temp_sda_s1_address -> temp_sda:address
	wire          mm_interconnect_2_temp_sda_s1_write;                                                       // mm_interconnect_2:temp_sda_s1_write -> temp_sda:write_n
	wire   [31:0] mm_interconnect_2_temp_sda_s1_writedata;                                                   // mm_interconnect_2:temp_sda_s1_writedata -> temp_sda:writedata
	wire          mm_interconnect_2_m2_ddr2_i2c_sda_s1_chipselect;                                           // mm_interconnect_2:m2_ddr2_i2c_sda_s1_chipselect -> m2_ddr2_i2c_sda:chipselect
	wire   [31:0] mm_interconnect_2_m2_ddr2_i2c_sda_s1_readdata;                                             // m2_ddr2_i2c_sda:readdata -> mm_interconnect_2:m2_ddr2_i2c_sda_s1_readdata
	wire    [1:0] mm_interconnect_2_m2_ddr2_i2c_sda_s1_address;                                              // mm_interconnect_2:m2_ddr2_i2c_sda_s1_address -> m2_ddr2_i2c_sda:address
	wire          mm_interconnect_2_m2_ddr2_i2c_sda_s1_write;                                                // mm_interconnect_2:m2_ddr2_i2c_sda_s1_write -> m2_ddr2_i2c_sda:write_n
	wire   [31:0] mm_interconnect_2_m2_ddr2_i2c_sda_s1_writedata;                                            // mm_interconnect_2:m2_ddr2_i2c_sda_s1_writedata -> m2_ddr2_i2c_sda:writedata
	wire          mm_interconnect_2_m2_ddr2_i2c_scl_s1_chipselect;                                           // mm_interconnect_2:m2_ddr2_i2c_scl_s1_chipselect -> m2_ddr2_i2c_scl:chipselect
	wire   [31:0] mm_interconnect_2_m2_ddr2_i2c_scl_s1_readdata;                                             // m2_ddr2_i2c_scl:readdata -> mm_interconnect_2:m2_ddr2_i2c_scl_s1_readdata
	wire    [1:0] mm_interconnect_2_m2_ddr2_i2c_scl_s1_address;                                              // mm_interconnect_2:m2_ddr2_i2c_scl_s1_address -> m2_ddr2_i2c_scl:address
	wire          mm_interconnect_2_m2_ddr2_i2c_scl_s1_write;                                                // mm_interconnect_2:m2_ddr2_i2c_scl_s1_write -> m2_ddr2_i2c_scl:write_n
	wire   [31:0] mm_interconnect_2_m2_ddr2_i2c_scl_s1_writedata;                                            // mm_interconnect_2:m2_ddr2_i2c_scl_s1_writedata -> m2_ddr2_i2c_scl:writedata
	wire   [31:0] mm_interconnect_2_csense_sdo_s1_readdata;                                                  // csense_sdo:readdata -> mm_interconnect_2:csense_sdo_s1_readdata
	wire    [1:0] mm_interconnect_2_csense_sdo_s1_address;                                                   // mm_interconnect_2:csense_sdo_s1_address -> csense_sdo:address
	wire          mm_interconnect_2_csense_sdi_s1_chipselect;                                                // mm_interconnect_2:csense_sdi_s1_chipselect -> csense_sdi:chipselect
	wire   [31:0] mm_interconnect_2_csense_sdi_s1_readdata;                                                  // csense_sdi:readdata -> mm_interconnect_2:csense_sdi_s1_readdata
	wire    [1:0] mm_interconnect_2_csense_sdi_s1_address;                                                   // mm_interconnect_2:csense_sdi_s1_address -> csense_sdi:address
	wire          mm_interconnect_2_csense_sdi_s1_write;                                                     // mm_interconnect_2:csense_sdi_s1_write -> csense_sdi:write_n
	wire   [31:0] mm_interconnect_2_csense_sdi_s1_writedata;                                                 // mm_interconnect_2:csense_sdi_s1_writedata -> csense_sdi:writedata
	wire          mm_interconnect_2_csense_sck_s1_chipselect;                                                // mm_interconnect_2:csense_sck_s1_chipselect -> csense_sck:chipselect
	wire   [31:0] mm_interconnect_2_csense_sck_s1_readdata;                                                  // csense_sck:readdata -> mm_interconnect_2:csense_sck_s1_readdata
	wire    [1:0] mm_interconnect_2_csense_sck_s1_address;                                                   // mm_interconnect_2:csense_sck_s1_address -> csense_sck:address
	wire          mm_interconnect_2_csense_sck_s1_write;                                                     // mm_interconnect_2:csense_sck_s1_write -> csense_sck:write_n
	wire   [31:0] mm_interconnect_2_csense_sck_s1_writedata;                                                 // mm_interconnect_2:csense_sck_s1_writedata -> csense_sck:writedata
	wire          mm_interconnect_2_csense_cs_n_s1_chipselect;                                               // mm_interconnect_2:csense_cs_n_s1_chipselect -> csense_cs_n:chipselect
	wire   [31:0] mm_interconnect_2_csense_cs_n_s1_readdata;                                                 // csense_cs_n:readdata -> mm_interconnect_2:csense_cs_n_s1_readdata
	wire    [1:0] mm_interconnect_2_csense_cs_n_s1_address;                                                  // mm_interconnect_2:csense_cs_n_s1_address -> csense_cs_n:address
	wire          mm_interconnect_2_csense_cs_n_s1_write;                                                    // mm_interconnect_2:csense_cs_n_s1_write -> csense_cs_n:write_n
	wire   [31:0] mm_interconnect_2_csense_cs_n_s1_writedata;                                                // mm_interconnect_2:csense_cs_n_s1_writedata -> csense_cs_n:writedata
	wire          mm_interconnect_2_csense_adc_fo_s1_chipselect;                                             // mm_interconnect_2:csense_adc_fo_s1_chipselect -> csense_adc_fo:chipselect
	wire   [31:0] mm_interconnect_2_csense_adc_fo_s1_readdata;                                               // csense_adc_fo:readdata -> mm_interconnect_2:csense_adc_fo_s1_readdata
	wire    [1:0] mm_interconnect_2_csense_adc_fo_s1_address;                                                // mm_interconnect_2:csense_adc_fo_s1_address -> csense_adc_fo:address
	wire          mm_interconnect_2_csense_adc_fo_s1_write;                                                  // mm_interconnect_2:csense_adc_fo_s1_write -> csense_adc_fo:write_n
	wire   [31:0] mm_interconnect_2_csense_adc_fo_s1_writedata;                                              // mm_interconnect_2:csense_adc_fo_s1_writedata -> csense_adc_fo:writedata
	wire          mm_interconnect_2_pio_led_painel_s1_chipselect;                                            // mm_interconnect_2:pio_LED_painel_s1_chipselect -> pio_LED_painel:chipselect
	wire   [31:0] mm_interconnect_2_pio_led_painel_s1_readdata;                                              // pio_LED_painel:readdata -> mm_interconnect_2:pio_LED_painel_s1_readdata
	wire    [1:0] mm_interconnect_2_pio_led_painel_s1_address;                                               // mm_interconnect_2:pio_LED_painel_s1_address -> pio_LED_painel:address
	wire          mm_interconnect_2_pio_led_painel_s1_write;                                                 // mm_interconnect_2:pio_LED_painel_s1_write -> pio_LED_painel:write_n
	wire   [31:0] mm_interconnect_2_pio_led_painel_s1_writedata;                                             // mm_interconnect_2:pio_LED_painel_s1_writedata -> pio_LED_painel:writedata
	wire   [31:0] mm_interconnect_2_rtcc_alarm_s1_readdata;                                                  // rtcc_alarm:readdata -> mm_interconnect_2:rtcc_alarm_s1_readdata
	wire    [1:0] mm_interconnect_2_rtcc_alarm_s1_address;                                                   // mm_interconnect_2:rtcc_alarm_s1_address -> rtcc_alarm:address
	wire   [31:0] mm_interconnect_2_rtcc_sdo_s1_readdata;                                                    // rtcc_sdo:readdata -> mm_interconnect_2:rtcc_sdo_s1_readdata
	wire    [1:0] mm_interconnect_2_rtcc_sdo_s1_address;                                                     // mm_interconnect_2:rtcc_sdo_s1_address -> rtcc_sdo:address
	wire          mm_interconnect_2_rtcc_sdi_s1_chipselect;                                                  // mm_interconnect_2:rtcc_sdi_s1_chipselect -> rtcc_sdi:chipselect
	wire   [31:0] mm_interconnect_2_rtcc_sdi_s1_readdata;                                                    // rtcc_sdi:readdata -> mm_interconnect_2:rtcc_sdi_s1_readdata
	wire    [1:0] mm_interconnect_2_rtcc_sdi_s1_address;                                                     // mm_interconnect_2:rtcc_sdi_s1_address -> rtcc_sdi:address
	wire          mm_interconnect_2_rtcc_sdi_s1_write;                                                       // mm_interconnect_2:rtcc_sdi_s1_write -> rtcc_sdi:write_n
	wire   [31:0] mm_interconnect_2_rtcc_sdi_s1_writedata;                                                   // mm_interconnect_2:rtcc_sdi_s1_writedata -> rtcc_sdi:writedata
	wire          mm_interconnect_2_rtcc_sck_s1_chipselect;                                                  // mm_interconnect_2:rtcc_sck_s1_chipselect -> rtcc_sck:chipselect
	wire   [31:0] mm_interconnect_2_rtcc_sck_s1_readdata;                                                    // rtcc_sck:readdata -> mm_interconnect_2:rtcc_sck_s1_readdata
	wire    [1:0] mm_interconnect_2_rtcc_sck_s1_address;                                                     // mm_interconnect_2:rtcc_sck_s1_address -> rtcc_sck:address
	wire          mm_interconnect_2_rtcc_sck_s1_write;                                                       // mm_interconnect_2:rtcc_sck_s1_write -> rtcc_sck:write_n
	wire   [31:0] mm_interconnect_2_rtcc_sck_s1_writedata;                                                   // mm_interconnect_2:rtcc_sck_s1_writedata -> rtcc_sck:writedata
	wire          mm_interconnect_2_rtcc_cs_n_s1_chipselect;                                                 // mm_interconnect_2:rtcc_cs_n_s1_chipselect -> rtcc_cs_n:chipselect
	wire   [31:0] mm_interconnect_2_rtcc_cs_n_s1_readdata;                                                   // rtcc_cs_n:readdata -> mm_interconnect_2:rtcc_cs_n_s1_readdata
	wire    [1:0] mm_interconnect_2_rtcc_cs_n_s1_address;                                                    // mm_interconnect_2:rtcc_cs_n_s1_address -> rtcc_cs_n:address
	wire          mm_interconnect_2_rtcc_cs_n_s1_write;                                                      // mm_interconnect_2:rtcc_cs_n_s1_write -> rtcc_cs_n:write_n
	wire   [31:0] mm_interconnect_2_rtcc_cs_n_s1_writedata;                                                  // mm_interconnect_2:rtcc_cs_n_s1_writedata -> rtcc_cs_n:writedata
	wire          mm_interconnect_2_rs232_uart_s1_chipselect;                                                // mm_interconnect_2:rs232_uart_s1_chipselect -> rs232_uart:chipselect
	wire   [15:0] mm_interconnect_2_rs232_uart_s1_readdata;                                                  // rs232_uart:readdata -> mm_interconnect_2:rs232_uart_s1_readdata
	wire    [2:0] mm_interconnect_2_rs232_uart_s1_address;                                                   // mm_interconnect_2:rs232_uart_s1_address -> rs232_uart:address
	wire          mm_interconnect_2_rs232_uart_s1_read;                                                      // mm_interconnect_2:rs232_uart_s1_read -> rs232_uart:read_n
	wire          mm_interconnect_2_rs232_uart_s1_begintransfer;                                             // mm_interconnect_2:rs232_uart_s1_begintransfer -> rs232_uart:begintransfer
	wire          mm_interconnect_2_rs232_uart_s1_write;                                                     // mm_interconnect_2:rs232_uart_s1_write -> rs232_uart:write_n
	wire   [15:0] mm_interconnect_2_rs232_uart_s1_writedata;                                                 // mm_interconnect_2:rs232_uart_s1_writedata -> rs232_uart:writedata
	wire          mm_interconnect_2_pio_ctrl_io_lvds_s1_chipselect;                                          // mm_interconnect_2:pio_ctrl_io_lvds_s1_chipselect -> pio_ctrl_io_lvds:chipselect
	wire   [31:0] mm_interconnect_2_pio_ctrl_io_lvds_s1_readdata;                                            // pio_ctrl_io_lvds:readdata -> mm_interconnect_2:pio_ctrl_io_lvds_s1_readdata
	wire    [1:0] mm_interconnect_2_pio_ctrl_io_lvds_s1_address;                                             // mm_interconnect_2:pio_ctrl_io_lvds_s1_address -> pio_ctrl_io_lvds:address
	wire          mm_interconnect_2_pio_ctrl_io_lvds_s1_write;                                               // mm_interconnect_2:pio_ctrl_io_lvds_s1_write -> pio_ctrl_io_lvds:write_n
	wire   [31:0] mm_interconnect_2_pio_ctrl_io_lvds_s1_writedata;                                           // mm_interconnect_2:pio_ctrl_io_lvds_s1_writedata -> pio_ctrl_io_lvds:writedata
	wire          m1_clock_bridge_m0_waitrequest;                                                            // mm_interconnect_3:m1_clock_bridge_m0_waitrequest -> m1_clock_bridge:m0_waitrequest
	wire  [255:0] m1_clock_bridge_m0_readdata;                                                               // mm_interconnect_3:m1_clock_bridge_m0_readdata -> m1_clock_bridge:m0_readdata
	wire          m1_clock_bridge_m0_debugaccess;                                                            // m1_clock_bridge:m0_debugaccess -> mm_interconnect_3:m1_clock_bridge_m0_debugaccess
	wire   [30:0] m1_clock_bridge_m0_address;                                                                // m1_clock_bridge:m0_address -> mm_interconnect_3:m1_clock_bridge_m0_address
	wire          m1_clock_bridge_m0_read;                                                                   // m1_clock_bridge:m0_read -> mm_interconnect_3:m1_clock_bridge_m0_read
	wire   [31:0] m1_clock_bridge_m0_byteenable;                                                             // m1_clock_bridge:m0_byteenable -> mm_interconnect_3:m1_clock_bridge_m0_byteenable
	wire          m1_clock_bridge_m0_readdatavalid;                                                          // mm_interconnect_3:m1_clock_bridge_m0_readdatavalid -> m1_clock_bridge:m0_readdatavalid
	wire  [255:0] m1_clock_bridge_m0_writedata;                                                              // m1_clock_bridge:m0_writedata -> mm_interconnect_3:m1_clock_bridge_m0_writedata
	wire          m1_clock_bridge_m0_write;                                                                  // m1_clock_bridge:m0_write -> mm_interconnect_3:m1_clock_bridge_m0_write
	wire    [2:0] m1_clock_bridge_m0_burstcount;                                                             // m1_clock_bridge:m0_burstcount -> mm_interconnect_3:m1_clock_bridge_m0_burstcount
	wire          mm_interconnect_3_m1_ddr2_memory_avl_beginbursttransfer;                                   // mm_interconnect_3:m1_ddr2_memory_avl_beginbursttransfer -> m1_ddr2_memory:avl_burstbegin
	wire  [255:0] mm_interconnect_3_m1_ddr2_memory_avl_readdata;                                             // m1_ddr2_memory:avl_rdata -> mm_interconnect_3:m1_ddr2_memory_avl_readdata
	wire          mm_interconnect_3_m1_ddr2_memory_avl_waitrequest;                                          // m1_ddr2_memory:avl_ready -> mm_interconnect_3:m1_ddr2_memory_avl_waitrequest
	wire   [25:0] mm_interconnect_3_m1_ddr2_memory_avl_address;                                              // mm_interconnect_3:m1_ddr2_memory_avl_address -> m1_ddr2_memory:avl_addr
	wire          mm_interconnect_3_m1_ddr2_memory_avl_read;                                                 // mm_interconnect_3:m1_ddr2_memory_avl_read -> m1_ddr2_memory:avl_read_req
	wire   [31:0] mm_interconnect_3_m1_ddr2_memory_avl_byteenable;                                           // mm_interconnect_3:m1_ddr2_memory_avl_byteenable -> m1_ddr2_memory:avl_be
	wire          mm_interconnect_3_m1_ddr2_memory_avl_readdatavalid;                                        // m1_ddr2_memory:avl_rdata_valid -> mm_interconnect_3:m1_ddr2_memory_avl_readdatavalid
	wire          mm_interconnect_3_m1_ddr2_memory_avl_write;                                                // mm_interconnect_3:m1_ddr2_memory_avl_write -> m1_ddr2_memory:avl_write_req
	wire  [255:0] mm_interconnect_3_m1_ddr2_memory_avl_writedata;                                            // mm_interconnect_3:m1_ddr2_memory_avl_writedata -> m1_ddr2_memory:avl_wdata
	wire    [7:0] mm_interconnect_3_m1_ddr2_memory_avl_burstcount;                                           // mm_interconnect_3:m1_ddr2_memory_avl_burstcount -> m1_ddr2_memory:avl_size
	wire          m1_ddr2_memory_afi_clk_clk;                                                                // m1_ddr2_memory:afi_clk -> [mm_interconnect_3:m1_ddr2_memory_afi_clk_clk, rst_controller_026:clk]
	wire          irq_mapper_receiver0_irq;                                                                  // COMM_Pedreiro_v1_01_1:buffers_interrupt_sender_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                  // COMM_Pedreiro_v1_01_2:buffers_interrupt_sender_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                  // COMM_Pedreiro_v1_01_3:buffers_interrupt_sender_irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                  // COMM_Pedreiro_v1_01_4:buffers_interrupt_sender_irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                                  // COMM_Pedreiro_v1_01_5:buffers_interrupt_sender_irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                                                  // COMM_Pedreiro_v1_01_6:buffers_interrupt_sender_irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                                                  // FTDI_USB3_0:ftdi_rx_interrupt_sender_irq -> irq_mapper:receiver6_irq
	wire          irq_mapper_receiver7_irq;                                                                  // FTDI_USB3_0:ftdi_tx_interrupt_sender_irq -> irq_mapper:receiver7_irq
	wire          irq_mapper_receiver8_irq;                                                                  // jtag_uart_0:av_irq -> irq_mapper:receiver8_irq
	wire          irq_mapper_receiver13_irq;                                                                 // COMM_Pedreiro_v1_01_1:rmap_interrupt_sender_irq -> irq_mapper:receiver13_irq
	wire          irq_mapper_receiver14_irq;                                                                 // COMM_Pedreiro_v1_01_2:rmap_interrupt_sender_irq -> irq_mapper:receiver14_irq
	wire          irq_mapper_receiver15_irq;                                                                 // COMM_Pedreiro_v1_01_3:rmap_interrupt_sender_irq -> irq_mapper:receiver15_irq
	wire          irq_mapper_receiver16_irq;                                                                 // COMM_Pedreiro_v1_01_4:rmap_interrupt_sender_irq -> irq_mapper:receiver16_irq
	wire          irq_mapper_receiver17_irq;                                                                 // COMM_Pedreiro_v1_01_5:rmap_interrupt_sender_irq -> irq_mapper:receiver17_irq
	wire          irq_mapper_receiver18_irq;                                                                 // COMM_Pedreiro_v1_01_6:rmap_interrupt_sender_irq -> irq_mapper:receiver18_irq
	wire   [31:0] nios2_gen2_0_irq_irq;                                                                      // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire          irq_mapper_receiver9_irq;                                                                  // irq_synchronizer:sender_irq -> irq_mapper:receiver9_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                             // timer_1ms:irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver10_irq;                                                                 // irq_synchronizer_001:sender_irq -> irq_mapper:receiver10_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                                                         // timer_1us:irq -> irq_synchronizer_001:receiver_irq
	wire          irq_mapper_receiver11_irq;                                                                 // irq_synchronizer_002:sender_irq -> irq_mapper:receiver11_irq
	wire    [0:0] irq_synchronizer_002_receiver_irq;                                                         // rs232_uart:irq -> irq_synchronizer_002:receiver_irq
	wire          irq_mapper_receiver12_irq;                                                                 // irq_synchronizer_003:sender_irq -> irq_mapper:receiver12_irq
	wire    [0:0] irq_synchronizer_003_receiver_irq;                                                         // sync:pre_sync_interrupt_sender_irq_o -> irq_synchronizer_003:receiver_irq
	wire          irq_mapper_receiver19_irq;                                                                 // irq_synchronizer_004:sender_irq -> irq_mapper:receiver19_irq
	wire    [0:0] irq_synchronizer_004_receiver_irq;                                                         // sync:sync_interrupt_sender_irq_o -> irq_synchronizer_004:receiver_irq
	wire          rst_controller_001_reset_out_reset;                                                        // rst_controller_001:reset_out -> [Altera_UP_SD_Card_Avalon_Interface_0:i_reset_n, mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_reset_source_sd_card_reset;                                                 // rst_controller:reset_source_sd_card_reset -> rst_controller_001:reset_in1
	wire          rst_controller_002_reset_out_reset;                                                        // rst_controller_002:reset_out -> [COMM_Pedreiro_v1_01_1:reset_sink_reset, mm_interconnect_0:COMM_Pedreiro_v1_01_1_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:rmap_mem_nfee_comm_1_reset_sink_reset_bridge_in_reset_reset, rmap_mem_nfee_comm_1:reset_i]
	wire          rst_controller_reset_source_comm_ch1_reset;                                                // rst_controller:reset_source_comm_ch1_reset -> [rst_controller_002:reset_in1, rst_controller_009:reset_in1, rst_controller_010:reset_in1]
	wire          rst_controller_003_reset_out_reset;                                                        // rst_controller_003:reset_out -> [COMM_Pedreiro_v1_01_2:reset_sink_reset, mm_interconnect_0:COMM_Pedreiro_v1_01_2_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:rmap_mem_nfee_comm_2_reset_sink_reset_bridge_in_reset_reset, rmap_mem_nfee_comm_2:reset_i]
	wire          rst_controller_reset_source_comm_ch2_reset;                                                // rst_controller:reset_source_comm_ch2_reset -> [rst_controller_003:reset_in1, rst_controller_009:reset_in2, rst_controller_011:reset_in1]
	wire          rst_controller_004_reset_out_reset;                                                        // rst_controller_004:reset_out -> [COMM_Pedreiro_v1_01_3:reset_sink_reset, mm_interconnect_0:COMM_Pedreiro_v1_01_3_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:rmap_mem_nfee_comm_3_reset_sink_reset_bridge_in_reset_reset, rmap_mem_nfee_comm_3:reset_i]
	wire          rst_controller_reset_source_comm_ch3_reset;                                                // rst_controller:reset_source_comm_ch3_reset -> [rst_controller_004:reset_in1, rst_controller_009:reset_in3, rst_controller_012:reset_in1]
	wire          rst_controller_005_reset_out_reset;                                                        // rst_controller_005:reset_out -> [COMM_Pedreiro_v1_01_4:reset_sink_reset, mm_interconnect_0:COMM_Pedreiro_v1_01_4_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:rmap_mem_nfee_comm_4_reset_sink_reset_bridge_in_reset_reset, rmap_mem_nfee_comm_4:reset_i]
	wire          rst_controller_reset_source_comm_ch4_reset;                                                // rst_controller:reset_source_comm_ch4_reset -> [rst_controller_005:reset_in1, rst_controller_009:reset_in4, rst_controller_013:reset_in1]
	wire          rst_controller_006_reset_out_reset;                                                        // rst_controller_006:reset_out -> [COMM_Pedreiro_v1_01_5:reset_sink_reset, mm_interconnect_0:COMM_Pedreiro_v1_01_5_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:rmap_mem_nfee_comm_5_reset_sink_reset_bridge_in_reset_reset, rmap_mem_nfee_comm_5:reset_i]
	wire          rst_controller_reset_source_comm_ch5_reset;                                                // rst_controller:reset_source_comm_ch5_reset -> [rst_controller_006:reset_in1, rst_controller_009:reset_in5, rst_controller_014:reset_in1]
	wire          rst_controller_007_reset_out_reset;                                                        // rst_controller_007:reset_out -> [COMM_Pedreiro_v1_01_6:reset_sink_reset, mm_interconnect_0:COMM_Pedreiro_v1_01_6_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:rmap_mem_nfee_comm_6_reset_sink_reset_bridge_in_reset_reset, rmap_mem_nfee_comm_6:reset_i]
	wire          rst_controller_reset_source_comm_ch6_reset;                                                // rst_controller:reset_source_comm_ch6_reset -> [rst_controller_007:reset_in1, rst_controller_009:reset_in6, rst_controller_015:reset_in1]
	wire          rst_controller_008_reset_out_reset;                                                        // rst_controller_008:reset_out -> [FTDI_USB3_0:reset_sink_reset, clock_bridge_afi_50:s0_reset, ddr2_address_span_extender:reset, jtag_uart_0:rst_n, m1_clock_bridge:s0_reset, mm_interconnect_0:FTDI_USB3_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_0:m1_clock_bridge_s0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:jtag_uart_0_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_translator:in_reset, sysid_qsys:reset_n]
	wire          rst_controller_008_reset_out_reset_req;                                                    // rst_controller_008:reset_req -> [onchip_memory:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_009_reset_out_reset;                                                        // rst_controller_009:reset_out -> RMAP_Echoing_0:reset_i
	wire          rst_controller_reset_source_comm_ch7_reset;                                                // rst_controller:reset_source_comm_ch7_reset -> [rst_controller_009:reset_in7, rst_controller_016:reset_in1, rst_controller_018:reset_in1]
	wire          rst_controller_reset_source_comm_ch8_reset;                                                // rst_controller:reset_source_comm_ch8_reset -> [rst_controller_009:reset_in8, rst_controller_017:reset_in1]
	wire          rst_controller_010_reset_out_reset;                                                        // rst_controller_010:reset_out -> SpaceWire_Channel_A:reset_i
	wire          rst_controller_011_reset_out_reset;                                                        // rst_controller_011:reset_out -> SpaceWire_Channel_B:reset_i
	wire          rst_controller_012_reset_out_reset;                                                        // rst_controller_012:reset_out -> SpaceWire_Channel_C:reset_i
	wire          rst_controller_013_reset_out_reset;                                                        // rst_controller_013:reset_out -> SpaceWire_Channel_D:reset_i
	wire          rst_controller_014_reset_out_reset;                                                        // rst_controller_014:reset_out -> SpaceWire_Channel_E:reset_i
	wire          rst_controller_015_reset_out_reset;                                                        // rst_controller_015:reset_out -> SpaceWire_Channel_F:reset_i
	wire          rst_controller_016_reset_out_reset;                                                        // rst_controller_016:reset_out -> SpaceWire_Channel_G:reset_i
	wire          rst_controller_017_reset_out_reset;                                                        // rst_controller_017:reset_out -> SpaceWire_Channel_H:reset_i
	wire          rst_controller_018_reset_out_reset;                                                        // rst_controller_018:reset_out -> SpaceWire_Glutton_0:reset_i
	wire          rst_controller_019_reset_out_reset;                                                        // rst_controller_019:reset_out -> [clock_bridge_afi_50:m0_reset, csense_adc_fo:reset_n, csense_cs_n:reset_n, csense_sck:reset_n, csense_sdi:reset_n, csense_sdo:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, m1_ddr2_i2c_scl:reset_n, m1_ddr2_i2c_sda:reset_n, m2_ddr2_i2c_scl:reset_n, m2_ddr2_i2c_sda:reset_n, mm_interconnect_2:clock_bridge_afi_50_m0_reset_reset_bridge_in_reset_reset, pio_BUTTON:reset_n, pio_DIP:reset_n, pio_EXT:reset_n, pio_LED:reset_n, pio_LED_painel:reset_n, pio_ctrl_io_lvds:reset_n, rst_controller:reset_sink_reset, rtcc_alarm:reset_n, rtcc_cs_n:reset_n, rtcc_sck:reset_n, rtcc_sdi:reset_n, rtcc_sdo:reset_n, sd_card_wp_n:reset_n, temp_scl:reset_n, temp_sda:reset_n, timer_1ms:reset_n, timer_1us:reset_n]
	wire          rst_controller_020_reset_out_reset;                                                        // rst_controller_020:reset_out -> [ext_flash:reset_reset, mm_interconnect_1:ext_flash_reset_reset_bridge_in_reset_reset, tristate_conduit_bridge_0:reset]
	wire          rst_controller_021_reset_out_reset;                                                        // rst_controller_021:reset_out -> [m1_clock_bridge:m0_reset, mm_interconnect_3:m1_clock_bridge_m0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_022_reset_out_reset;                                                        // rst_controller_022:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, mm_interconnect_1:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator_001:in_reset]
	wire          rst_controller_022_reset_out_reset_req;                                                    // rst_controller_022:reset_req -> [nios2_gen2_0:reset_req, rst_translator_001:reset_req_in]
	wire          rst_controller_023_reset_out_reset;                                                        // rst_controller_023:reset_out -> [irq_synchronizer_002:receiver_reset, mm_interconnect_2:rs232_uart_reset_reset_bridge_in_reset_reset, rs232_uart:reset_n]
	wire          rst_controller_reset_source_rs232_reset;                                                   // rst_controller:reset_source_rs232_reset -> rst_controller_023:reset_in1
	wire          rst_controller_024_reset_out_reset;                                                        // rst_controller_024:reset_out -> [irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, mm_interconnect_2:sync_reset_reset_bridge_in_reset_reset, sync:reset_sink_reset_i]
	wire          rst_controller_reset_source_sync_reset;                                                    // rst_controller:reset_source_sync_reset -> rst_controller_024:reset_in1
	wire          rst_controller_025_reset_out_reset;                                                        // rst_controller_025:reset_out -> [mm_interconnect_0:m2_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:m2_ddr2_memory_soft_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_026_reset_out_reset;                                                        // rst_controller_026:reset_out -> [mm_interconnect_3:m1_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_3:m1_ddr2_memory_soft_reset_reset_bridge_in_reset_reset]

	Altera_UP_SD_Card_Avalon_Interface altera_up_sd_card_avalon_interface_0 (
		.i_avalon_chip_select (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address),     //                    .address
		.i_avalon_read        (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read),        //                    .read
		.i_avalon_write       (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write),       //                    .write
		.i_avalon_byteenable  (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable),  //                    .byteenable
		.i_avalon_writedata   (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata),   //                    .writedata
		.o_avalon_readdata    (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata),    //                    .readdata
		.o_avalon_waitrequest (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest), //                    .waitrequest
		.i_clock              (clk50_clk),                                                                              //                 clk.clk
		.i_reset_n            (~rst_controller_001_reset_out_reset),                                                    //               reset.reset_n
		.b_SD_cmd             (sd_card_ip_b_SD_cmd),                                                                    //         conduit_end.export
		.b_SD_dat             (sd_card_ip_b_SD_dat),                                                                    //                    .export
		.b_SD_dat3            (sd_card_ip_b_SD_dat3),                                                                   //                    .export
		.o_SD_clock           (sd_card_ip_o_SD_clock)                                                                   //                    .export
	);

	comm_v1_80_top comm_pedreiro_v1_01_1 (
		.reset_sink_reset                     (rst_controller_002_reset_out_reset),                                                        //                        reset_sink.reset
		.sync_channel                         (comm_a_sync_end_sync_channel_signal),                                                       //                  sync_conduit_end.sync_channel_signal
		.rmap_interrupt_sender_irq            (irq_mapper_receiver13_irq),                                                                 //             rmap_interrupt_sender.irq
		.buffers_interrupt_sender_irq         (irq_mapper_receiver0_irq),                                                                  //          buffers_interrupt_sender.irq
		.clock_sink_100_clk                   (m2_ddr2_memory_afi_half_clk_clk),                                                           //                    clock_sink_100.clk
		.clock_sink_200_clk                   (m2_ddr2_memory_afi_clk_clk),                                                                //                    clock_sink_200.clk
		.avalon_slave_windowing_address       (mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_address),                    //            avalon_slave_windowing.address
		.avalon_slave_windowing_write         (mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_write),                      //                                  .write
		.avalon_slave_windowing_read          (mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_read),                       //                                  .read
		.avalon_slave_windowing_writedata     (mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_writedata),                  //                                  .writedata
		.avalon_slave_windowing_byteenable    (mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_byteenable),                 //                                  .byteenable
		.avalon_slave_windowing_readdata      (mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_readdata),                   //                                  .readdata
		.avalon_slave_windowing_waitrequest   (mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_waitrequest),                //                                  .waitrequest
		.avm_left_buffer_readdata_i           (comm_pedreiro_v1_01_1_avalon_mm_left_buffer_master_readdata),                               //      avalon_mm_left_buffer_master.readdata
		.avm_left_buffer_waitrequest_i        (comm_pedreiro_v1_01_1_avalon_mm_left_buffer_master_waitrequest),                            //                                  .waitrequest
		.avm_left_buffer_address_o            (comm_pedreiro_v1_01_1_avalon_mm_left_buffer_master_address),                                //                                  .address
		.avm_left_buffer_read_o               (comm_pedreiro_v1_01_1_avalon_mm_left_buffer_master_read),                                   //                                  .read
		.avm_right_buffer_readdata_i          (comm_pedreiro_v1_01_1_avalon_mm_right_buffer_master_readdata),                              //     avalon_mm_right_buffer_master.readdata
		.avm_right_buffer_waitrequest_i       (comm_pedreiro_v1_01_1_avalon_mm_right_buffer_master_waitrequest),                           //                                  .waitrequest
		.avm_right_buffer_address_o           (comm_pedreiro_v1_01_1_avalon_mm_right_buffer_master_address),                               //                                  .address
		.avm_right_buffer_read_o              (comm_pedreiro_v1_01_1_avalon_mm_right_buffer_master_read),                                  //                                  .read
		.spw_link_status_started_i            (spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_started_signal),          //  conduit_end_spacewire_controller.spw_link_status_started_signal
		.spw_link_status_connecting_i         (spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_connecting_signal),       //                                  .spw_link_status_connecting_signal
		.spw_link_status_running_i            (spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_running_signal),          //                                  .spw_link_status_running_signal
		.spw_link_error_errdisc_i             (spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),           //                                  .spw_link_error_errdisc_signal
		.spw_link_error_errpar_i              (spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errpar_signal),            //                                  .spw_link_error_errpar_signal
		.spw_link_error_erresc_i              (spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_erresc_signal),            //                                  .spw_link_error_erresc_signal
		.spw_link_error_errcred_i             (spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errcred_signal),           //                                  .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_i           (spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),         //                                  .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_i           (spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),         //                                  .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_i           (spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),         //                                  .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_i         (spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),       //                                  .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_i         (spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),       //                                  .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_i          (spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),        //                                  .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_i          (spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),        //                                  .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_i           (spacewire_channel_a_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),         //                                  .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_i         (spacewire_channel_a_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal),       //                                  .spw_data_tx_status_txhalff_signal
		.spw_link_command_autostart_o         (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_link_command_autostart_signal),  //                                  .spw_link_command_autostart_signal
		.spw_link_command_linkstart_o         (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),  //                                  .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_o           (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),    //                                  .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_o          (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),   //                                  .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_o            (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),     //                                  .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_o            (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),     //                                  .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_o            (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),     //                                  .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_o         (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),  //                                  .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_o        (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal), //                                  .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_o         (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),  //                                  .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_o         (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal),  //                                  .spw_data_tx_command_txdata_signal
		.measurements_channel                 (comm_a_measurements_conduit_end_measurements_channel_signal),                               //          measurements_conduit_end.measurements_channel_signal
		.fee_rmap_echo_en_o                   (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_echo_en_signal),                        //     conduit_end_fee_rmap_echo_out.echo_en_signal
		.fee_rmap_echo_id_en_o                (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_echo_id_en_signal),                     //                                  .echo_id_en_signal
		.fee_rmap_incoming_fifo_wrdata_flag_o (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal),      //                                  .incoming_fifo_wrdata_flag_signal
		.fee_rmap_incoming_fifo_wrdata_data_o (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal),      //                                  .incoming_fifo_wrdata_data_signal
		.fee_rmap_incoming_fifo_wrreq_o       (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal),            //                                  .incoming_fifo_wrreq_signal
		.fee_rmap_outgoing_fifo_wrdata_flag_o (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal),      //                                  .outgoing_fifo_wrdata_flag_signal
		.fee_rmap_outgoing_fifo_wrdata_data_o (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal),      //                                  .outgoing_fifo_wrdata_data_signal
		.fee_rmap_outgoing_fifo_wrreq_o       (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal),            //                                  .outgoing_fifo_wrreq_signal
		.fee_codec_rmap_wr_waitrequest_i      (rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal),                   // conduit_end_fee_rmap_master_codec.wr_waitrequest_signal
		.fee_codec_rmap_readdata_i            (rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_readdata_signal),                         //                                  .readdata_signal
		.fee_codec_rmap_rd_waitrequest_i      (rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal),                   //                                  .rd_waitrequest_signal
		.fee_codec_rmap_wr_address_o          (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_wr_address_signal),                 //                                  .wr_address_signal
		.fee_codec_rmap_write_o               (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_write_signal),                      //                                  .write_signal
		.fee_codec_rmap_writedata_o           (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_writedata_signal),                  //                                  .writedata_signal
		.fee_codec_rmap_rd_address_o          (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_rd_address_signal),                 //                                  .rd_address_signal
		.fee_codec_rmap_read_o                (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_read_signal),                       //                                  .read_signal
		.fee_hk_rmap_wr_waitrequest_i         (rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal),                   //    conduit_end_fee_rmap_master_hk.wr_waitrequest_signal
		.fee_hk_rmap_readdata_i               (rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_readdata_signal),                         //                                  .readdata_signal
		.fee_hk_rmap_rd_waitrequest_i         (rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal),                   //                                  .rd_waitrequest_signal
		.fee_hk_rmap_wr_address_o             (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_wr_address_signal),                    //                                  .wr_address_signal
		.fee_hk_rmap_write_o                  (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_write_signal),                         //                                  .write_signal
		.fee_hk_rmap_writedata_o              (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_writedata_signal),                     //                                  .writedata_signal
		.fee_hk_rmap_rd_address_o             (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_rd_address_signal),                    //                                  .rd_address_signal
		.fee_hk_rmap_read_o                   (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_read_signal),                          //                                  .read_signal
		.channel_hk_timecode_control_o        (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_timecode_control_signal),                  //        conduit_end_channel_hk_out.timecode_control_signal
		.channel_hk_timecode_time_o           (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_timecode_time_signal),                     //                                  .timecode_time_signal
		.channel_hk_rmap_target_status_o      (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_rmap_target_status_signal),                //                                  .rmap_target_status_signal
		.channel_hk_rmap_target_indicate_o    (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_rmap_target_indicate_signal),              //                                  .rmap_target_indicate_signal
		.channel_hk_spw_link_escape_err_o     (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_escape_err_signal),               //                                  .spw_link_escape_err_signal
		.channel_hk_spw_link_credit_err_o     (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_credit_err_signal),               //                                  .spw_link_credit_err_signal
		.channel_hk_spw_link_parity_err_o     (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_parity_err_signal),               //                                  .spw_link_parity_err_signal
		.channel_hk_spw_link_disconnect_o     (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_disconnect_signal),               //                                  .spw_link_disconnect_signal
		.channel_hk_spw_link_running_o        (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_running_signal),                  //                                  .spw_link_running_signal
		.channel_hk_frame_counter_o           (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_frame_counter_signal),                     //                                  .frame_counter_signal
		.channel_hk_frame_number_o            (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_frame_number_signal),                      //                                  .frame_number_signal
		.channel_hk_err_win_wrong_x_coord_o   (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal),             //                                  .err_win_wrong_x_coord_signal
		.channel_hk_err_win_wrong_y_coord_o   (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal),             //                                  .err_win_wrong_y_coord_signal
		.channel_hk_err_e_side_buffer_full_o  (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_e_side_buffer_full_signal),            //                                  .err_e_side_buffer_full_signal
		.channel_hk_err_f_side_buffer_full_o  (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_f_side_buffer_full_signal),            //                                  .err_f_side_buffer_full_signal
		.channel_hk_err_invalid_ccd_mode_o    (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal),              //                                  .err_invalid_ccd_mode_signal
		.channel_win_mem_addr_offset_o        (comm_pedreiro_v1_01_1_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal)          //  conduit_end_rmap_avm_configs_out.win_mem_addr_offset_signal
	);

	comm_v1_80_top comm_pedreiro_v1_01_2 (
		.reset_sink_reset                     (rst_controller_003_reset_out_reset),                                                        //                        reset_sink.reset
		.sync_channel                         (comm_b_sync_end_sync_channel_signal),                                                       //                  sync_conduit_end.sync_channel_signal
		.rmap_interrupt_sender_irq            (irq_mapper_receiver14_irq),                                                                 //             rmap_interrupt_sender.irq
		.buffers_interrupt_sender_irq         (irq_mapper_receiver1_irq),                                                                  //          buffers_interrupt_sender.irq
		.clock_sink_100_clk                   (m2_ddr2_memory_afi_half_clk_clk),                                                           //                    clock_sink_100.clk
		.clock_sink_200_clk                   (m2_ddr2_memory_afi_clk_clk),                                                                //                    clock_sink_200.clk
		.avalon_slave_windowing_address       (mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_address),                    //            avalon_slave_windowing.address
		.avalon_slave_windowing_write         (mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_write),                      //                                  .write
		.avalon_slave_windowing_read          (mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_read),                       //                                  .read
		.avalon_slave_windowing_writedata     (mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_writedata),                  //                                  .writedata
		.avalon_slave_windowing_byteenable    (mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_byteenable),                 //                                  .byteenable
		.avalon_slave_windowing_readdata      (mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_readdata),                   //                                  .readdata
		.avalon_slave_windowing_waitrequest   (mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_waitrequest),                //                                  .waitrequest
		.avm_left_buffer_readdata_i           (comm_pedreiro_v1_01_2_avalon_mm_left_buffer_master_readdata),                               //      avalon_mm_left_buffer_master.readdata
		.avm_left_buffer_waitrequest_i        (comm_pedreiro_v1_01_2_avalon_mm_left_buffer_master_waitrequest),                            //                                  .waitrequest
		.avm_left_buffer_address_o            (comm_pedreiro_v1_01_2_avalon_mm_left_buffer_master_address),                                //                                  .address
		.avm_left_buffer_read_o               (comm_pedreiro_v1_01_2_avalon_mm_left_buffer_master_read),                                   //                                  .read
		.avm_right_buffer_readdata_i          (comm_pedreiro_v1_01_2_avalon_mm_right_buffer_master_readdata),                              //     avalon_mm_right_buffer_master.readdata
		.avm_right_buffer_waitrequest_i       (comm_pedreiro_v1_01_2_avalon_mm_right_buffer_master_waitrequest),                           //                                  .waitrequest
		.avm_right_buffer_address_o           (comm_pedreiro_v1_01_2_avalon_mm_right_buffer_master_address),                               //                                  .address
		.avm_right_buffer_read_o              (comm_pedreiro_v1_01_2_avalon_mm_right_buffer_master_read),                                  //                                  .read
		.spw_link_status_started_i            (spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_started_signal),          //  conduit_end_spacewire_controller.spw_link_status_started_signal
		.spw_link_status_connecting_i         (spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_connecting_signal),       //                                  .spw_link_status_connecting_signal
		.spw_link_status_running_i            (spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_running_signal),          //                                  .spw_link_status_running_signal
		.spw_link_error_errdisc_i             (spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),           //                                  .spw_link_error_errdisc_signal
		.spw_link_error_errpar_i              (spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errpar_signal),            //                                  .spw_link_error_errpar_signal
		.spw_link_error_erresc_i              (spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_erresc_signal),            //                                  .spw_link_error_erresc_signal
		.spw_link_error_errcred_i             (spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errcred_signal),           //                                  .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_i           (spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),         //                                  .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_i           (spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),         //                                  .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_i           (spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),         //                                  .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_i         (spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),       //                                  .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_i         (spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),       //                                  .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_i          (spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),        //                                  .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_i          (spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),        //                                  .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_i           (spacewire_channel_b_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),         //                                  .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_i         (spacewire_channel_b_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal),       //                                  .spw_data_tx_status_txhalff_signal
		.spw_link_command_autostart_o         (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_link_command_autostart_signal),  //                                  .spw_link_command_autostart_signal
		.spw_link_command_linkstart_o         (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),  //                                  .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_o           (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),    //                                  .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_o          (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),   //                                  .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_o            (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),     //                                  .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_o            (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),     //                                  .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_o            (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),     //                                  .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_o         (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),  //                                  .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_o        (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal), //                                  .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_o         (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),  //                                  .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_o         (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal),  //                                  .spw_data_tx_command_txdata_signal
		.measurements_channel                 (comm_b_measurements_conduit_end_measurements_channel_signal),                               //          measurements_conduit_end.measurements_channel_signal
		.fee_rmap_echo_en_o                   (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_echo_en_signal),                        //     conduit_end_fee_rmap_echo_out.echo_en_signal
		.fee_rmap_echo_id_en_o                (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_echo_id_en_signal),                     //                                  .echo_id_en_signal
		.fee_rmap_incoming_fifo_wrdata_flag_o (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal),      //                                  .incoming_fifo_wrdata_flag_signal
		.fee_rmap_incoming_fifo_wrdata_data_o (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal),      //                                  .incoming_fifo_wrdata_data_signal
		.fee_rmap_incoming_fifo_wrreq_o       (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal),            //                                  .incoming_fifo_wrreq_signal
		.fee_rmap_outgoing_fifo_wrdata_flag_o (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal),      //                                  .outgoing_fifo_wrdata_flag_signal
		.fee_rmap_outgoing_fifo_wrdata_data_o (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal),      //                                  .outgoing_fifo_wrdata_data_signal
		.fee_rmap_outgoing_fifo_wrreq_o       (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal),            //                                  .outgoing_fifo_wrreq_signal
		.fee_codec_rmap_wr_waitrequest_i      (rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal),                   // conduit_end_fee_rmap_master_codec.wr_waitrequest_signal
		.fee_codec_rmap_readdata_i            (rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_readdata_signal),                         //                                  .readdata_signal
		.fee_codec_rmap_rd_waitrequest_i      (rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal),                   //                                  .rd_waitrequest_signal
		.fee_codec_rmap_wr_address_o          (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_wr_address_signal),                 //                                  .wr_address_signal
		.fee_codec_rmap_write_o               (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_write_signal),                      //                                  .write_signal
		.fee_codec_rmap_writedata_o           (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_writedata_signal),                  //                                  .writedata_signal
		.fee_codec_rmap_rd_address_o          (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_rd_address_signal),                 //                                  .rd_address_signal
		.fee_codec_rmap_read_o                (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_read_signal),                       //                                  .read_signal
		.fee_hk_rmap_wr_waitrequest_i         (rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal),                   //    conduit_end_fee_rmap_master_hk.wr_waitrequest_signal
		.fee_hk_rmap_readdata_i               (rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_readdata_signal),                         //                                  .readdata_signal
		.fee_hk_rmap_rd_waitrequest_i         (rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal),                   //                                  .rd_waitrequest_signal
		.fee_hk_rmap_wr_address_o             (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_wr_address_signal),                    //                                  .wr_address_signal
		.fee_hk_rmap_write_o                  (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_write_signal),                         //                                  .write_signal
		.fee_hk_rmap_writedata_o              (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_writedata_signal),                     //                                  .writedata_signal
		.fee_hk_rmap_rd_address_o             (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_rd_address_signal),                    //                                  .rd_address_signal
		.fee_hk_rmap_read_o                   (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_read_signal),                          //                                  .read_signal
		.channel_hk_timecode_control_o        (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_timecode_control_signal),                  //        conduit_end_channel_hk_out.timecode_control_signal
		.channel_hk_timecode_time_o           (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_timecode_time_signal),                     //                                  .timecode_time_signal
		.channel_hk_rmap_target_status_o      (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_rmap_target_status_signal),                //                                  .rmap_target_status_signal
		.channel_hk_rmap_target_indicate_o    (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_rmap_target_indicate_signal),              //                                  .rmap_target_indicate_signal
		.channel_hk_spw_link_escape_err_o     (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_escape_err_signal),               //                                  .spw_link_escape_err_signal
		.channel_hk_spw_link_credit_err_o     (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_credit_err_signal),               //                                  .spw_link_credit_err_signal
		.channel_hk_spw_link_parity_err_o     (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_parity_err_signal),               //                                  .spw_link_parity_err_signal
		.channel_hk_spw_link_disconnect_o     (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_disconnect_signal),               //                                  .spw_link_disconnect_signal
		.channel_hk_spw_link_running_o        (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_running_signal),                  //                                  .spw_link_running_signal
		.channel_hk_frame_counter_o           (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_frame_counter_signal),                     //                                  .frame_counter_signal
		.channel_hk_frame_number_o            (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_frame_number_signal),                      //                                  .frame_number_signal
		.channel_hk_err_win_wrong_x_coord_o   (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal),             //                                  .err_win_wrong_x_coord_signal
		.channel_hk_err_win_wrong_y_coord_o   (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal),             //                                  .err_win_wrong_y_coord_signal
		.channel_hk_err_e_side_buffer_full_o  (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_e_side_buffer_full_signal),            //                                  .err_e_side_buffer_full_signal
		.channel_hk_err_f_side_buffer_full_o  (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_f_side_buffer_full_signal),            //                                  .err_f_side_buffer_full_signal
		.channel_hk_err_invalid_ccd_mode_o    (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal),              //                                  .err_invalid_ccd_mode_signal
		.channel_win_mem_addr_offset_o        (comm_pedreiro_v1_01_2_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal)          //  conduit_end_rmap_avm_configs_out.win_mem_addr_offset_signal
	);

	comm_v1_80_top comm_pedreiro_v1_01_3 (
		.reset_sink_reset                     (rst_controller_004_reset_out_reset),                                                        //                        reset_sink.reset
		.sync_channel                         (comm_c_sync_end_sync_channel_signal),                                                       //                  sync_conduit_end.sync_channel_signal
		.rmap_interrupt_sender_irq            (irq_mapper_receiver15_irq),                                                                 //             rmap_interrupt_sender.irq
		.buffers_interrupt_sender_irq         (irq_mapper_receiver2_irq),                                                                  //          buffers_interrupt_sender.irq
		.clock_sink_100_clk                   (m2_ddr2_memory_afi_half_clk_clk),                                                           //                    clock_sink_100.clk
		.clock_sink_200_clk                   (m2_ddr2_memory_afi_clk_clk),                                                                //                    clock_sink_200.clk
		.avalon_slave_windowing_address       (mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_address),                    //            avalon_slave_windowing.address
		.avalon_slave_windowing_write         (mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_write),                      //                                  .write
		.avalon_slave_windowing_read          (mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_read),                       //                                  .read
		.avalon_slave_windowing_writedata     (mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_writedata),                  //                                  .writedata
		.avalon_slave_windowing_byteenable    (mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_byteenable),                 //                                  .byteenable
		.avalon_slave_windowing_readdata      (mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_readdata),                   //                                  .readdata
		.avalon_slave_windowing_waitrequest   (mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_waitrequest),                //                                  .waitrequest
		.avm_left_buffer_readdata_i           (comm_pedreiro_v1_01_3_avalon_mm_left_buffer_master_readdata),                               //      avalon_mm_left_buffer_master.readdata
		.avm_left_buffer_waitrequest_i        (comm_pedreiro_v1_01_3_avalon_mm_left_buffer_master_waitrequest),                            //                                  .waitrequest
		.avm_left_buffer_address_o            (comm_pedreiro_v1_01_3_avalon_mm_left_buffer_master_address),                                //                                  .address
		.avm_left_buffer_read_o               (comm_pedreiro_v1_01_3_avalon_mm_left_buffer_master_read),                                   //                                  .read
		.avm_right_buffer_readdata_i          (comm_pedreiro_v1_01_3_avalon_mm_right_buffer_master_readdata),                              //     avalon_mm_right_buffer_master.readdata
		.avm_right_buffer_waitrequest_i       (comm_pedreiro_v1_01_3_avalon_mm_right_buffer_master_waitrequest),                           //                                  .waitrequest
		.avm_right_buffer_address_o           (comm_pedreiro_v1_01_3_avalon_mm_right_buffer_master_address),                               //                                  .address
		.avm_right_buffer_read_o              (comm_pedreiro_v1_01_3_avalon_mm_right_buffer_master_read),                                  //                                  .read
		.spw_link_status_started_i            (spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_started_signal),          //  conduit_end_spacewire_controller.spw_link_status_started_signal
		.spw_link_status_connecting_i         (spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_connecting_signal),       //                                  .spw_link_status_connecting_signal
		.spw_link_status_running_i            (spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_running_signal),          //                                  .spw_link_status_running_signal
		.spw_link_error_errdisc_i             (spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),           //                                  .spw_link_error_errdisc_signal
		.spw_link_error_errpar_i              (spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errpar_signal),            //                                  .spw_link_error_errpar_signal
		.spw_link_error_erresc_i              (spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_erresc_signal),            //                                  .spw_link_error_erresc_signal
		.spw_link_error_errcred_i             (spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errcred_signal),           //                                  .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_i           (spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),         //                                  .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_i           (spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),         //                                  .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_i           (spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),         //                                  .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_i         (spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),       //                                  .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_i         (spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),       //                                  .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_i          (spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),        //                                  .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_i          (spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),        //                                  .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_i           (spacewire_channel_c_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),         //                                  .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_i         (spacewire_channel_c_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal),       //                                  .spw_data_tx_status_txhalff_signal
		.spw_link_command_autostart_o         (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_link_command_autostart_signal),  //                                  .spw_link_command_autostart_signal
		.spw_link_command_linkstart_o         (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),  //                                  .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_o           (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),    //                                  .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_o          (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),   //                                  .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_o            (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),     //                                  .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_o            (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),     //                                  .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_o            (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),     //                                  .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_o         (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),  //                                  .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_o        (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal), //                                  .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_o         (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),  //                                  .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_o         (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal),  //                                  .spw_data_tx_command_txdata_signal
		.measurements_channel                 (comm_c_measurements_conduit_end_measurements_channel_signal),                               //          measurements_conduit_end.measurements_channel_signal
		.fee_rmap_echo_en_o                   (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_echo_en_signal),                        //     conduit_end_fee_rmap_echo_out.echo_en_signal
		.fee_rmap_echo_id_en_o                (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_echo_id_en_signal),                     //                                  .echo_id_en_signal
		.fee_rmap_incoming_fifo_wrdata_flag_o (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal),      //                                  .incoming_fifo_wrdata_flag_signal
		.fee_rmap_incoming_fifo_wrdata_data_o (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal),      //                                  .incoming_fifo_wrdata_data_signal
		.fee_rmap_incoming_fifo_wrreq_o       (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal),            //                                  .incoming_fifo_wrreq_signal
		.fee_rmap_outgoing_fifo_wrdata_flag_o (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal),      //                                  .outgoing_fifo_wrdata_flag_signal
		.fee_rmap_outgoing_fifo_wrdata_data_o (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal),      //                                  .outgoing_fifo_wrdata_data_signal
		.fee_rmap_outgoing_fifo_wrreq_o       (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal),            //                                  .outgoing_fifo_wrreq_signal
		.fee_codec_rmap_wr_waitrequest_i      (rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal),                   // conduit_end_fee_rmap_master_codec.wr_waitrequest_signal
		.fee_codec_rmap_readdata_i            (rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_readdata_signal),                         //                                  .readdata_signal
		.fee_codec_rmap_rd_waitrequest_i      (rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal),                   //                                  .rd_waitrequest_signal
		.fee_codec_rmap_wr_address_o          (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_wr_address_signal),                 //                                  .wr_address_signal
		.fee_codec_rmap_write_o               (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_write_signal),                      //                                  .write_signal
		.fee_codec_rmap_writedata_o           (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_writedata_signal),                  //                                  .writedata_signal
		.fee_codec_rmap_rd_address_o          (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_rd_address_signal),                 //                                  .rd_address_signal
		.fee_codec_rmap_read_o                (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_read_signal),                       //                                  .read_signal
		.fee_hk_rmap_wr_waitrequest_i         (rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal),                   //    conduit_end_fee_rmap_master_hk.wr_waitrequest_signal
		.fee_hk_rmap_readdata_i               (rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_readdata_signal),                         //                                  .readdata_signal
		.fee_hk_rmap_rd_waitrequest_i         (rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal),                   //                                  .rd_waitrequest_signal
		.fee_hk_rmap_wr_address_o             (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_wr_address_signal),                    //                                  .wr_address_signal
		.fee_hk_rmap_write_o                  (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_write_signal),                         //                                  .write_signal
		.fee_hk_rmap_writedata_o              (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_writedata_signal),                     //                                  .writedata_signal
		.fee_hk_rmap_rd_address_o             (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_rd_address_signal),                    //                                  .rd_address_signal
		.fee_hk_rmap_read_o                   (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_read_signal),                          //                                  .read_signal
		.channel_hk_timecode_control_o        (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_timecode_control_signal),                  //        conduit_end_channel_hk_out.timecode_control_signal
		.channel_hk_timecode_time_o           (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_timecode_time_signal),                     //                                  .timecode_time_signal
		.channel_hk_rmap_target_status_o      (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_rmap_target_status_signal),                //                                  .rmap_target_status_signal
		.channel_hk_rmap_target_indicate_o    (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_rmap_target_indicate_signal),              //                                  .rmap_target_indicate_signal
		.channel_hk_spw_link_escape_err_o     (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_escape_err_signal),               //                                  .spw_link_escape_err_signal
		.channel_hk_spw_link_credit_err_o     (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_credit_err_signal),               //                                  .spw_link_credit_err_signal
		.channel_hk_spw_link_parity_err_o     (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_parity_err_signal),               //                                  .spw_link_parity_err_signal
		.channel_hk_spw_link_disconnect_o     (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_disconnect_signal),               //                                  .spw_link_disconnect_signal
		.channel_hk_spw_link_running_o        (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_running_signal),                  //                                  .spw_link_running_signal
		.channel_hk_frame_counter_o           (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_frame_counter_signal),                     //                                  .frame_counter_signal
		.channel_hk_frame_number_o            (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_frame_number_signal),                      //                                  .frame_number_signal
		.channel_hk_err_win_wrong_x_coord_o   (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal),             //                                  .err_win_wrong_x_coord_signal
		.channel_hk_err_win_wrong_y_coord_o   (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal),             //                                  .err_win_wrong_y_coord_signal
		.channel_hk_err_e_side_buffer_full_o  (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_e_side_buffer_full_signal),            //                                  .err_e_side_buffer_full_signal
		.channel_hk_err_f_side_buffer_full_o  (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_f_side_buffer_full_signal),            //                                  .err_f_side_buffer_full_signal
		.channel_hk_err_invalid_ccd_mode_o    (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal),              //                                  .err_invalid_ccd_mode_signal
		.channel_win_mem_addr_offset_o        (comm_pedreiro_v1_01_3_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal)          //  conduit_end_rmap_avm_configs_out.win_mem_addr_offset_signal
	);

	comm_v1_80_top comm_pedreiro_v1_01_4 (
		.reset_sink_reset                     (rst_controller_005_reset_out_reset),                                                        //                        reset_sink.reset
		.sync_channel                         (comm_d_sync_end_sync_channel_signal),                                                       //                  sync_conduit_end.sync_channel_signal
		.rmap_interrupt_sender_irq            (irq_mapper_receiver16_irq),                                                                 //             rmap_interrupt_sender.irq
		.buffers_interrupt_sender_irq         (irq_mapper_receiver3_irq),                                                                  //          buffers_interrupt_sender.irq
		.clock_sink_100_clk                   (m2_ddr2_memory_afi_half_clk_clk),                                                           //                    clock_sink_100.clk
		.clock_sink_200_clk                   (m2_ddr2_memory_afi_clk_clk),                                                                //                    clock_sink_200.clk
		.avalon_slave_windowing_address       (mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_address),                    //            avalon_slave_windowing.address
		.avalon_slave_windowing_write         (mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_write),                      //                                  .write
		.avalon_slave_windowing_read          (mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_read),                       //                                  .read
		.avalon_slave_windowing_writedata     (mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_writedata),                  //                                  .writedata
		.avalon_slave_windowing_byteenable    (mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_byteenable),                 //                                  .byteenable
		.avalon_slave_windowing_readdata      (mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_readdata),                   //                                  .readdata
		.avalon_slave_windowing_waitrequest   (mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_waitrequest),                //                                  .waitrequest
		.avm_left_buffer_readdata_i           (comm_pedreiro_v1_01_4_avalon_mm_left_buffer_master_readdata),                               //      avalon_mm_left_buffer_master.readdata
		.avm_left_buffer_waitrequest_i        (comm_pedreiro_v1_01_4_avalon_mm_left_buffer_master_waitrequest),                            //                                  .waitrequest
		.avm_left_buffer_address_o            (comm_pedreiro_v1_01_4_avalon_mm_left_buffer_master_address),                                //                                  .address
		.avm_left_buffer_read_o               (comm_pedreiro_v1_01_4_avalon_mm_left_buffer_master_read),                                   //                                  .read
		.avm_right_buffer_readdata_i          (comm_pedreiro_v1_01_4_avalon_mm_right_buffer_master_readdata),                              //     avalon_mm_right_buffer_master.readdata
		.avm_right_buffer_waitrequest_i       (comm_pedreiro_v1_01_4_avalon_mm_right_buffer_master_waitrequest),                           //                                  .waitrequest
		.avm_right_buffer_address_o           (comm_pedreiro_v1_01_4_avalon_mm_right_buffer_master_address),                               //                                  .address
		.avm_right_buffer_read_o              (comm_pedreiro_v1_01_4_avalon_mm_right_buffer_master_read),                                  //                                  .read
		.spw_link_status_started_i            (spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_started_signal),          //  conduit_end_spacewire_controller.spw_link_status_started_signal
		.spw_link_status_connecting_i         (spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_connecting_signal),       //                                  .spw_link_status_connecting_signal
		.spw_link_status_running_i            (spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_running_signal),          //                                  .spw_link_status_running_signal
		.spw_link_error_errdisc_i             (spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),           //                                  .spw_link_error_errdisc_signal
		.spw_link_error_errpar_i              (spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errpar_signal),            //                                  .spw_link_error_errpar_signal
		.spw_link_error_erresc_i              (spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_erresc_signal),            //                                  .spw_link_error_erresc_signal
		.spw_link_error_errcred_i             (spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errcred_signal),           //                                  .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_i           (spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),         //                                  .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_i           (spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),         //                                  .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_i           (spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),         //                                  .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_i         (spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),       //                                  .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_i         (spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),       //                                  .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_i          (spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),        //                                  .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_i          (spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),        //                                  .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_i           (spacewire_channel_d_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),         //                                  .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_i         (spacewire_channel_d_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal),       //                                  .spw_data_tx_status_txhalff_signal
		.spw_link_command_autostart_o         (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_link_command_autostart_signal),  //                                  .spw_link_command_autostart_signal
		.spw_link_command_linkstart_o         (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),  //                                  .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_o           (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),    //                                  .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_o          (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),   //                                  .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_o            (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),     //                                  .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_o            (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),     //                                  .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_o            (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),     //                                  .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_o         (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),  //                                  .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_o        (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal), //                                  .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_o         (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),  //                                  .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_o         (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal),  //                                  .spw_data_tx_command_txdata_signal
		.measurements_channel                 (comm_d_measurements_conduit_end_measurements_channel_signal),                               //          measurements_conduit_end.measurements_channel_signal
		.fee_rmap_echo_en_o                   (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_echo_en_signal),                        //     conduit_end_fee_rmap_echo_out.echo_en_signal
		.fee_rmap_echo_id_en_o                (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_echo_id_en_signal),                     //                                  .echo_id_en_signal
		.fee_rmap_incoming_fifo_wrdata_flag_o (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal),      //                                  .incoming_fifo_wrdata_flag_signal
		.fee_rmap_incoming_fifo_wrdata_data_o (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal),      //                                  .incoming_fifo_wrdata_data_signal
		.fee_rmap_incoming_fifo_wrreq_o       (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal),            //                                  .incoming_fifo_wrreq_signal
		.fee_rmap_outgoing_fifo_wrdata_flag_o (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal),      //                                  .outgoing_fifo_wrdata_flag_signal
		.fee_rmap_outgoing_fifo_wrdata_data_o (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal),      //                                  .outgoing_fifo_wrdata_data_signal
		.fee_rmap_outgoing_fifo_wrreq_o       (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal),            //                                  .outgoing_fifo_wrreq_signal
		.fee_codec_rmap_wr_waitrequest_i      (rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal),                   // conduit_end_fee_rmap_master_codec.wr_waitrequest_signal
		.fee_codec_rmap_readdata_i            (rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_readdata_signal),                         //                                  .readdata_signal
		.fee_codec_rmap_rd_waitrequest_i      (rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal),                   //                                  .rd_waitrequest_signal
		.fee_codec_rmap_wr_address_o          (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_wr_address_signal),                 //                                  .wr_address_signal
		.fee_codec_rmap_write_o               (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_write_signal),                      //                                  .write_signal
		.fee_codec_rmap_writedata_o           (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_writedata_signal),                  //                                  .writedata_signal
		.fee_codec_rmap_rd_address_o          (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_rd_address_signal),                 //                                  .rd_address_signal
		.fee_codec_rmap_read_o                (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_read_signal),                       //                                  .read_signal
		.fee_hk_rmap_wr_waitrequest_i         (rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal),                   //    conduit_end_fee_rmap_master_hk.wr_waitrequest_signal
		.fee_hk_rmap_readdata_i               (rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_readdata_signal),                         //                                  .readdata_signal
		.fee_hk_rmap_rd_waitrequest_i         (rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal),                   //                                  .rd_waitrequest_signal
		.fee_hk_rmap_wr_address_o             (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_wr_address_signal),                    //                                  .wr_address_signal
		.fee_hk_rmap_write_o                  (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_write_signal),                         //                                  .write_signal
		.fee_hk_rmap_writedata_o              (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_writedata_signal),                     //                                  .writedata_signal
		.fee_hk_rmap_rd_address_o             (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_rd_address_signal),                    //                                  .rd_address_signal
		.fee_hk_rmap_read_o                   (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_read_signal),                          //                                  .read_signal
		.channel_hk_timecode_control_o        (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_timecode_control_signal),                  //        conduit_end_channel_hk_out.timecode_control_signal
		.channel_hk_timecode_time_o           (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_timecode_time_signal),                     //                                  .timecode_time_signal
		.channel_hk_rmap_target_status_o      (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_rmap_target_status_signal),                //                                  .rmap_target_status_signal
		.channel_hk_rmap_target_indicate_o    (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_rmap_target_indicate_signal),              //                                  .rmap_target_indicate_signal
		.channel_hk_spw_link_escape_err_o     (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_escape_err_signal),               //                                  .spw_link_escape_err_signal
		.channel_hk_spw_link_credit_err_o     (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_credit_err_signal),               //                                  .spw_link_credit_err_signal
		.channel_hk_spw_link_parity_err_o     (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_parity_err_signal),               //                                  .spw_link_parity_err_signal
		.channel_hk_spw_link_disconnect_o     (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_disconnect_signal),               //                                  .spw_link_disconnect_signal
		.channel_hk_spw_link_running_o        (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_running_signal),                  //                                  .spw_link_running_signal
		.channel_hk_frame_counter_o           (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_frame_counter_signal),                     //                                  .frame_counter_signal
		.channel_hk_frame_number_o            (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_frame_number_signal),                      //                                  .frame_number_signal
		.channel_hk_err_win_wrong_x_coord_o   (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal),             //                                  .err_win_wrong_x_coord_signal
		.channel_hk_err_win_wrong_y_coord_o   (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal),             //                                  .err_win_wrong_y_coord_signal
		.channel_hk_err_e_side_buffer_full_o  (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_e_side_buffer_full_signal),            //                                  .err_e_side_buffer_full_signal
		.channel_hk_err_f_side_buffer_full_o  (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_f_side_buffer_full_signal),            //                                  .err_f_side_buffer_full_signal
		.channel_hk_err_invalid_ccd_mode_o    (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal),              //                                  .err_invalid_ccd_mode_signal
		.channel_win_mem_addr_offset_o        (comm_pedreiro_v1_01_4_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal)          //  conduit_end_rmap_avm_configs_out.win_mem_addr_offset_signal
	);

	comm_v1_80_top comm_pedreiro_v1_01_5 (
		.reset_sink_reset                     (rst_controller_006_reset_out_reset),                                                        //                        reset_sink.reset
		.sync_channel                         (comm_e_sync_end_sync_channel_signal),                                                       //                  sync_conduit_end.sync_channel_signal
		.rmap_interrupt_sender_irq            (irq_mapper_receiver17_irq),                                                                 //             rmap_interrupt_sender.irq
		.buffers_interrupt_sender_irq         (irq_mapper_receiver4_irq),                                                                  //          buffers_interrupt_sender.irq
		.clock_sink_100_clk                   (m2_ddr2_memory_afi_half_clk_clk),                                                           //                    clock_sink_100.clk
		.clock_sink_200_clk                   (m2_ddr2_memory_afi_clk_clk),                                                                //                    clock_sink_200.clk
		.avalon_slave_windowing_address       (mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_address),                    //            avalon_slave_windowing.address
		.avalon_slave_windowing_write         (mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_write),                      //                                  .write
		.avalon_slave_windowing_read          (mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_read),                       //                                  .read
		.avalon_slave_windowing_writedata     (mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_writedata),                  //                                  .writedata
		.avalon_slave_windowing_byteenable    (mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_byteenable),                 //                                  .byteenable
		.avalon_slave_windowing_readdata      (mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_readdata),                   //                                  .readdata
		.avalon_slave_windowing_waitrequest   (mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_waitrequest),                //                                  .waitrequest
		.avm_left_buffer_readdata_i           (comm_pedreiro_v1_01_5_avalon_mm_left_buffer_master_readdata),                               //      avalon_mm_left_buffer_master.readdata
		.avm_left_buffer_waitrequest_i        (comm_pedreiro_v1_01_5_avalon_mm_left_buffer_master_waitrequest),                            //                                  .waitrequest
		.avm_left_buffer_address_o            (comm_pedreiro_v1_01_5_avalon_mm_left_buffer_master_address),                                //                                  .address
		.avm_left_buffer_read_o               (comm_pedreiro_v1_01_5_avalon_mm_left_buffer_master_read),                                   //                                  .read
		.avm_right_buffer_readdata_i          (comm_pedreiro_v1_01_5_avalon_mm_right_buffer_master_readdata),                              //     avalon_mm_right_buffer_master.readdata
		.avm_right_buffer_waitrequest_i       (comm_pedreiro_v1_01_5_avalon_mm_right_buffer_master_waitrequest),                           //                                  .waitrequest
		.avm_right_buffer_address_o           (comm_pedreiro_v1_01_5_avalon_mm_right_buffer_master_address),                               //                                  .address
		.avm_right_buffer_read_o              (comm_pedreiro_v1_01_5_avalon_mm_right_buffer_master_read),                                  //                                  .read
		.spw_link_status_started_i            (spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_started_signal),          //  conduit_end_spacewire_controller.spw_link_status_started_signal
		.spw_link_status_connecting_i         (spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_connecting_signal),       //                                  .spw_link_status_connecting_signal
		.spw_link_status_running_i            (spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_running_signal),          //                                  .spw_link_status_running_signal
		.spw_link_error_errdisc_i             (spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),           //                                  .spw_link_error_errdisc_signal
		.spw_link_error_errpar_i              (spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errpar_signal),            //                                  .spw_link_error_errpar_signal
		.spw_link_error_erresc_i              (spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_erresc_signal),            //                                  .spw_link_error_erresc_signal
		.spw_link_error_errcred_i             (spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errcred_signal),           //                                  .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_i           (spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),         //                                  .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_i           (spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),         //                                  .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_i           (spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),         //                                  .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_i         (spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),       //                                  .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_i         (spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),       //                                  .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_i          (spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),        //                                  .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_i          (spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),        //                                  .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_i           (spacewire_channel_e_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),         //                                  .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_i         (spacewire_channel_e_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal),       //                                  .spw_data_tx_status_txhalff_signal
		.spw_link_command_autostart_o         (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_link_command_autostart_signal),  //                                  .spw_link_command_autostart_signal
		.spw_link_command_linkstart_o         (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),  //                                  .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_o           (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),    //                                  .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_o          (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),   //                                  .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_o            (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),     //                                  .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_o            (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),     //                                  .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_o            (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),     //                                  .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_o         (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),  //                                  .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_o        (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal), //                                  .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_o         (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),  //                                  .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_o         (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal),  //                                  .spw_data_tx_command_txdata_signal
		.measurements_channel                 (comm_e_measurements_conduit_end_measurements_channel_signal),                               //          measurements_conduit_end.measurements_channel_signal
		.fee_rmap_echo_en_o                   (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_echo_en_signal),                        //     conduit_end_fee_rmap_echo_out.echo_en_signal
		.fee_rmap_echo_id_en_o                (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_echo_id_en_signal),                     //                                  .echo_id_en_signal
		.fee_rmap_incoming_fifo_wrdata_flag_o (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal),      //                                  .incoming_fifo_wrdata_flag_signal
		.fee_rmap_incoming_fifo_wrdata_data_o (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal),      //                                  .incoming_fifo_wrdata_data_signal
		.fee_rmap_incoming_fifo_wrreq_o       (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal),            //                                  .incoming_fifo_wrreq_signal
		.fee_rmap_outgoing_fifo_wrdata_flag_o (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal),      //                                  .outgoing_fifo_wrdata_flag_signal
		.fee_rmap_outgoing_fifo_wrdata_data_o (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal),      //                                  .outgoing_fifo_wrdata_data_signal
		.fee_rmap_outgoing_fifo_wrreq_o       (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal),            //                                  .outgoing_fifo_wrreq_signal
		.fee_codec_rmap_wr_waitrequest_i      (rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal),                   // conduit_end_fee_rmap_master_codec.wr_waitrequest_signal
		.fee_codec_rmap_readdata_i            (rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_readdata_signal),                         //                                  .readdata_signal
		.fee_codec_rmap_rd_waitrequest_i      (rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal),                   //                                  .rd_waitrequest_signal
		.fee_codec_rmap_wr_address_o          (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_wr_address_signal),                 //                                  .wr_address_signal
		.fee_codec_rmap_write_o               (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_write_signal),                      //                                  .write_signal
		.fee_codec_rmap_writedata_o           (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_writedata_signal),                  //                                  .writedata_signal
		.fee_codec_rmap_rd_address_o          (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_rd_address_signal),                 //                                  .rd_address_signal
		.fee_codec_rmap_read_o                (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_read_signal),                       //                                  .read_signal
		.fee_hk_rmap_wr_waitrequest_i         (rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal),                   //    conduit_end_fee_rmap_master_hk.wr_waitrequest_signal
		.fee_hk_rmap_readdata_i               (rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_readdata_signal),                         //                                  .readdata_signal
		.fee_hk_rmap_rd_waitrequest_i         (rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal),                   //                                  .rd_waitrequest_signal
		.fee_hk_rmap_wr_address_o             (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_wr_address_signal),                    //                                  .wr_address_signal
		.fee_hk_rmap_write_o                  (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_write_signal),                         //                                  .write_signal
		.fee_hk_rmap_writedata_o              (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_writedata_signal),                     //                                  .writedata_signal
		.fee_hk_rmap_rd_address_o             (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_rd_address_signal),                    //                                  .rd_address_signal
		.fee_hk_rmap_read_o                   (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_read_signal),                          //                                  .read_signal
		.channel_hk_timecode_control_o        (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_timecode_control_signal),                  //        conduit_end_channel_hk_out.timecode_control_signal
		.channel_hk_timecode_time_o           (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_timecode_time_signal),                     //                                  .timecode_time_signal
		.channel_hk_rmap_target_status_o      (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_rmap_target_status_signal),                //                                  .rmap_target_status_signal
		.channel_hk_rmap_target_indicate_o    (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_rmap_target_indicate_signal),              //                                  .rmap_target_indicate_signal
		.channel_hk_spw_link_escape_err_o     (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_escape_err_signal),               //                                  .spw_link_escape_err_signal
		.channel_hk_spw_link_credit_err_o     (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_credit_err_signal),               //                                  .spw_link_credit_err_signal
		.channel_hk_spw_link_parity_err_o     (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_parity_err_signal),               //                                  .spw_link_parity_err_signal
		.channel_hk_spw_link_disconnect_o     (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_disconnect_signal),               //                                  .spw_link_disconnect_signal
		.channel_hk_spw_link_running_o        (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_running_signal),                  //                                  .spw_link_running_signal
		.channel_hk_frame_counter_o           (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_frame_counter_signal),                     //                                  .frame_counter_signal
		.channel_hk_frame_number_o            (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_frame_number_signal),                      //                                  .frame_number_signal
		.channel_hk_err_win_wrong_x_coord_o   (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal),             //                                  .err_win_wrong_x_coord_signal
		.channel_hk_err_win_wrong_y_coord_o   (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal),             //                                  .err_win_wrong_y_coord_signal
		.channel_hk_err_e_side_buffer_full_o  (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_e_side_buffer_full_signal),            //                                  .err_e_side_buffer_full_signal
		.channel_hk_err_f_side_buffer_full_o  (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_f_side_buffer_full_signal),            //                                  .err_f_side_buffer_full_signal
		.channel_hk_err_invalid_ccd_mode_o    (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal),              //                                  .err_invalid_ccd_mode_signal
		.channel_win_mem_addr_offset_o        (comm_pedreiro_v1_01_5_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal)          //  conduit_end_rmap_avm_configs_out.win_mem_addr_offset_signal
	);

	comm_v1_80_top comm_pedreiro_v1_01_6 (
		.reset_sink_reset                     (rst_controller_007_reset_out_reset),                                                        //                        reset_sink.reset
		.sync_channel                         (comm_f_sync_end_sync_channel_signal),                                                       //                  sync_conduit_end.sync_channel_signal
		.rmap_interrupt_sender_irq            (irq_mapper_receiver18_irq),                                                                 //             rmap_interrupt_sender.irq
		.buffers_interrupt_sender_irq         (irq_mapper_receiver5_irq),                                                                  //          buffers_interrupt_sender.irq
		.clock_sink_100_clk                   (m2_ddr2_memory_afi_half_clk_clk),                                                           //                    clock_sink_100.clk
		.clock_sink_200_clk                   (m2_ddr2_memory_afi_clk_clk),                                                                //                    clock_sink_200.clk
		.avalon_slave_windowing_address       (mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_address),                    //            avalon_slave_windowing.address
		.avalon_slave_windowing_write         (mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_write),                      //                                  .write
		.avalon_slave_windowing_read          (mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_read),                       //                                  .read
		.avalon_slave_windowing_writedata     (mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_writedata),                  //                                  .writedata
		.avalon_slave_windowing_byteenable    (mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_byteenable),                 //                                  .byteenable
		.avalon_slave_windowing_readdata      (mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_readdata),                   //                                  .readdata
		.avalon_slave_windowing_waitrequest   (mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_waitrequest),                //                                  .waitrequest
		.avm_left_buffer_readdata_i           (comm_pedreiro_v1_01_6_avalon_mm_left_buffer_master_readdata),                               //      avalon_mm_left_buffer_master.readdata
		.avm_left_buffer_waitrequest_i        (comm_pedreiro_v1_01_6_avalon_mm_left_buffer_master_waitrequest),                            //                                  .waitrequest
		.avm_left_buffer_address_o            (comm_pedreiro_v1_01_6_avalon_mm_left_buffer_master_address),                                //                                  .address
		.avm_left_buffer_read_o               (comm_pedreiro_v1_01_6_avalon_mm_left_buffer_master_read),                                   //                                  .read
		.avm_right_buffer_readdata_i          (comm_pedreiro_v1_01_6_avalon_mm_right_buffer_master_readdata),                              //     avalon_mm_right_buffer_master.readdata
		.avm_right_buffer_waitrequest_i       (comm_pedreiro_v1_01_6_avalon_mm_right_buffer_master_waitrequest),                           //                                  .waitrequest
		.avm_right_buffer_address_o           (comm_pedreiro_v1_01_6_avalon_mm_right_buffer_master_address),                               //                                  .address
		.avm_right_buffer_read_o              (comm_pedreiro_v1_01_6_avalon_mm_right_buffer_master_read),                                  //                                  .read
		.spw_link_status_started_i            (spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_started_signal),          //  conduit_end_spacewire_controller.spw_link_status_started_signal
		.spw_link_status_connecting_i         (spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_connecting_signal),       //                                  .spw_link_status_connecting_signal
		.spw_link_status_running_i            (spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_running_signal),          //                                  .spw_link_status_running_signal
		.spw_link_error_errdisc_i             (spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),           //                                  .spw_link_error_errdisc_signal
		.spw_link_error_errpar_i              (spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errpar_signal),            //                                  .spw_link_error_errpar_signal
		.spw_link_error_erresc_i              (spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_erresc_signal),            //                                  .spw_link_error_erresc_signal
		.spw_link_error_errcred_i             (spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errcred_signal),           //                                  .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_i           (spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),         //                                  .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_i           (spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),         //                                  .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_i           (spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),         //                                  .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_i         (spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),       //                                  .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_i         (spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),       //                                  .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_i          (spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),        //                                  .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_i          (spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),        //                                  .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_i           (spacewire_channel_f_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),         //                                  .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_i         (spacewire_channel_f_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal),       //                                  .spw_data_tx_status_txhalff_signal
		.spw_link_command_autostart_o         (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_link_command_autostart_signal),  //                                  .spw_link_command_autostart_signal
		.spw_link_command_linkstart_o         (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),  //                                  .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_o           (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),    //                                  .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_o          (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),   //                                  .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_o            (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),     //                                  .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_o            (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),     //                                  .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_o            (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),     //                                  .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_o         (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),  //                                  .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_o        (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal), //                                  .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_o         (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),  //                                  .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_o         (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal),  //                                  .spw_data_tx_command_txdata_signal
		.measurements_channel                 (comm_f_measurements_conduit_end_measurements_channel_signal),                               //          measurements_conduit_end.measurements_channel_signal
		.fee_rmap_echo_en_o                   (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_echo_en_signal),                        //     conduit_end_fee_rmap_echo_out.echo_en_signal
		.fee_rmap_echo_id_en_o                (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_echo_id_en_signal),                     //                                  .echo_id_en_signal
		.fee_rmap_incoming_fifo_wrdata_flag_o (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal),      //                                  .incoming_fifo_wrdata_flag_signal
		.fee_rmap_incoming_fifo_wrdata_data_o (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal),      //                                  .incoming_fifo_wrdata_data_signal
		.fee_rmap_incoming_fifo_wrreq_o       (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal),            //                                  .incoming_fifo_wrreq_signal
		.fee_rmap_outgoing_fifo_wrdata_flag_o (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal),      //                                  .outgoing_fifo_wrdata_flag_signal
		.fee_rmap_outgoing_fifo_wrdata_data_o (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal),      //                                  .outgoing_fifo_wrdata_data_signal
		.fee_rmap_outgoing_fifo_wrreq_o       (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal),            //                                  .outgoing_fifo_wrreq_signal
		.fee_codec_rmap_wr_waitrequest_i      (rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal),                   // conduit_end_fee_rmap_master_codec.wr_waitrequest_signal
		.fee_codec_rmap_readdata_i            (rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_readdata_signal),                         //                                  .readdata_signal
		.fee_codec_rmap_rd_waitrequest_i      (rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal),                   //                                  .rd_waitrequest_signal
		.fee_codec_rmap_wr_address_o          (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_wr_address_signal),                 //                                  .wr_address_signal
		.fee_codec_rmap_write_o               (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_write_signal),                      //                                  .write_signal
		.fee_codec_rmap_writedata_o           (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_writedata_signal),                  //                                  .writedata_signal
		.fee_codec_rmap_rd_address_o          (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_rd_address_signal),                 //                                  .rd_address_signal
		.fee_codec_rmap_read_o                (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_read_signal),                       //                                  .read_signal
		.fee_hk_rmap_wr_waitrequest_i         (rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal),                   //    conduit_end_fee_rmap_master_hk.wr_waitrequest_signal
		.fee_hk_rmap_readdata_i               (rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_readdata_signal),                         //                                  .readdata_signal
		.fee_hk_rmap_rd_waitrequest_i         (rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal),                   //                                  .rd_waitrequest_signal
		.fee_hk_rmap_wr_address_o             (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_wr_address_signal),                    //                                  .wr_address_signal
		.fee_hk_rmap_write_o                  (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_write_signal),                         //                                  .write_signal
		.fee_hk_rmap_writedata_o              (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_writedata_signal),                     //                                  .writedata_signal
		.fee_hk_rmap_rd_address_o             (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_rd_address_signal),                    //                                  .rd_address_signal
		.fee_hk_rmap_read_o                   (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_read_signal),                          //                                  .read_signal
		.channel_hk_timecode_control_o        (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_timecode_control_signal),                  //        conduit_end_channel_hk_out.timecode_control_signal
		.channel_hk_timecode_time_o           (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_timecode_time_signal),                     //                                  .timecode_time_signal
		.channel_hk_rmap_target_status_o      (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_rmap_target_status_signal),                //                                  .rmap_target_status_signal
		.channel_hk_rmap_target_indicate_o    (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_rmap_target_indicate_signal),              //                                  .rmap_target_indicate_signal
		.channel_hk_spw_link_escape_err_o     (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_escape_err_signal),               //                                  .spw_link_escape_err_signal
		.channel_hk_spw_link_credit_err_o     (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_credit_err_signal),               //                                  .spw_link_credit_err_signal
		.channel_hk_spw_link_parity_err_o     (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_parity_err_signal),               //                                  .spw_link_parity_err_signal
		.channel_hk_spw_link_disconnect_o     (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_disconnect_signal),               //                                  .spw_link_disconnect_signal
		.channel_hk_spw_link_running_o        (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_running_signal),                  //                                  .spw_link_running_signal
		.channel_hk_frame_counter_o           (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_frame_counter_signal),                     //                                  .frame_counter_signal
		.channel_hk_frame_number_o            (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_frame_number_signal),                      //                                  .frame_number_signal
		.channel_hk_err_win_wrong_x_coord_o   (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal),             //                                  .err_win_wrong_x_coord_signal
		.channel_hk_err_win_wrong_y_coord_o   (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal),             //                                  .err_win_wrong_y_coord_signal
		.channel_hk_err_e_side_buffer_full_o  (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_e_side_buffer_full_signal),            //                                  .err_e_side_buffer_full_signal
		.channel_hk_err_f_side_buffer_full_o  (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_f_side_buffer_full_signal),            //                                  .err_f_side_buffer_full_signal
		.channel_hk_err_invalid_ccd_mode_o    (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal),              //                                  .err_invalid_ccd_mode_signal
		.channel_win_mem_addr_offset_o        (comm_pedreiro_v1_01_6_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal)          //  conduit_end_rmap_avm_configs_out.win_mem_addr_offset_signal
	);

	ftdi_usb3_top ftdi_usb3_0 (
		.clock_sink_clk                  (m2_ddr2_memory_afi_half_clk_clk),                               //               clock_sink.clk
		.ftdi_clock_sink_clk             (ftdi_clk_clk),                                                  //          ftdi_clock_sink.clk
		.reset_sink_reset                (rst_controller_008_reset_out_reset),                            //               reset_sink.reset
		.umft_data_bus                   (umft601a_pins_umft_data_signal),                                //        conduit_umft_pins.umft_data_signal
		.umft_reset_n_pin                (umft601a_pins_umft_reset_n_signal),                             //                         .umft_reset_n_signal
		.umft_rxf_n_pin                  (umft601a_pins_umft_rxf_n_signal),                               //                         .umft_rxf_n_signal
		.umft_clock_pin                  (umft601a_pins_umft_clock_signal),                               //                         .umft_clock_signal
		.umft_wakeup_n_pin               (umft601a_pins_umft_wakeup_n_signal),                            //                         .umft_wakeup_n_signal
		.umft_be_bus                     (umft601a_pins_umft_be_signal),                                  //                         .umft_be_signal
		.umft_txe_n_pin                  (umft601a_pins_umft_txe_n_signal),                               //                         .umft_txe_n_signal
		.umft_gpio_bus                   (umft601a_pins_umft_gpio_bus_signal),                            //                         .umft_gpio_bus_signal
		.umft_wr_n_pin                   (umft601a_pins_umft_wr_n_signal),                                //                         .umft_wr_n_signal
		.umft_rd_n_pin                   (umft601a_pins_umft_rd_n_signal),                                //                         .umft_rd_n_signal
		.umft_oe_n_pin                   (umft601a_pins_umft_oe_n_signal),                                //                         .umft_oe_n_signal
		.umft_siwu_n_pin                 (umft601a_pins_umft_siwu_n_signal),                              //                         .umft_siwu_n_signal
		.avalon_slave_config_address     (mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_address),     //      avalon_slave_config.address
		.avalon_slave_config_byteenable  (mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_byteenable),  //                         .byteenable
		.avalon_slave_config_write       (mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_write),       //                         .write
		.avalon_slave_config_writedata   (mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_writedata),   //                         .writedata
		.avalon_slave_config_read        (mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_read),        //                         .read
		.avalon_slave_config_readdata    (mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_readdata),    //                         .readdata
		.avalon_slave_config_waitrequest (mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_waitrequest), //                         .waitrequest
		.avalon_master_data_readdata     (ftdi_usb3_0_avalon_master_data_readdata),                       //       avalon_master_data.readdata
		.avalon_master_data_waitrequest  (ftdi_usb3_0_avalon_master_data_waitrequest),                    //                         .waitrequest
		.avalon_master_data_address      (ftdi_usb3_0_avalon_master_data_address),                        //                         .address
		.avalon_master_data_read         (ftdi_usb3_0_avalon_master_data_read),                           //                         .read
		.avalon_master_data_write        (ftdi_usb3_0_avalon_master_data_write),                          //                         .write
		.avalon_master_data_writedata    (ftdi_usb3_0_avalon_master_data_writedata),                      //                         .writedata
		.ftdi_rx_interrupt_sender_irq    (irq_mapper_receiver6_irq),                                      // ftdi_rx_interrupt_sender.irq
		.ftdi_tx_interrupt_sender_irq    (irq_mapper_receiver7_irq)                                       // ftdi_tx_interrupt_sender.irq
	);

	rmpe_rmap_echoing_top rmap_echoing_0 (
		.reset_i                                (rst_controller_009_reset_out_reset),                                                   //                       reset_sink.reset
		.clk_100_i                              (m2_ddr2_memory_afi_half_clk_clk),                                                      //                clock_sink_100mhz.clk
		.fee_0_rmap_echo_en_i                   (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_echo_en_signal),                   //   conduit_end_fee_0_rmap_echo_in.echo_en_signal
		.fee_0_rmap_echo_id_en_i                (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_echo_id_en_signal),                //                                 .echo_id_en_signal
		.fee_0_rmap_incoming_fifo_wrdata_flag_i (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal), //                                 .incoming_fifo_wrdata_flag_signal
		.fee_0_rmap_incoming_fifo_wrdata_data_i (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal), //                                 .incoming_fifo_wrdata_data_signal
		.fee_0_rmap_incoming_fifo_wrreq_i       (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal),       //                                 .incoming_fifo_wrreq_signal
		.fee_0_rmap_outgoing_fifo_wrdata_flag_i (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal), //                                 .outgoing_fifo_wrdata_flag_signal
		.fee_0_rmap_outgoing_fifo_wrdata_data_i (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal), //                                 .outgoing_fifo_wrdata_data_signal
		.fee_0_rmap_outgoing_fifo_wrreq_i       (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal),       //                                 .outgoing_fifo_wrreq_signal
		.fee_1_rmap_echo_en_i                   (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_echo_en_signal),                   //   conduit_end_fee_1_rmap_echo_in.echo_en_signal
		.fee_1_rmap_echo_id_en_i                (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_echo_id_en_signal),                //                                 .echo_id_en_signal
		.fee_1_rmap_incoming_fifo_wrdata_flag_i (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal), //                                 .incoming_fifo_wrdata_flag_signal
		.fee_1_rmap_incoming_fifo_wrdata_data_i (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal), //                                 .incoming_fifo_wrdata_data_signal
		.fee_1_rmap_incoming_fifo_wrreq_i       (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal),       //                                 .incoming_fifo_wrreq_signal
		.fee_1_rmap_outgoing_fifo_wrdata_flag_i (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal), //                                 .outgoing_fifo_wrdata_flag_signal
		.fee_1_rmap_outgoing_fifo_wrdata_data_i (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal), //                                 .outgoing_fifo_wrdata_data_signal
		.fee_1_rmap_outgoing_fifo_wrreq_i       (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal),       //                                 .outgoing_fifo_wrreq_signal
		.fee_2_rmap_echo_en_i                   (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_echo_en_signal),                   //   conduit_end_fee_2_rmap_echo_in.echo_en_signal
		.fee_2_rmap_echo_id_en_i                (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_echo_id_en_signal),                //                                 .echo_id_en_signal
		.fee_2_rmap_incoming_fifo_wrdata_flag_i (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal), //                                 .incoming_fifo_wrdata_flag_signal
		.fee_2_rmap_incoming_fifo_wrdata_data_i (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal), //                                 .incoming_fifo_wrdata_data_signal
		.fee_2_rmap_incoming_fifo_wrreq_i       (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal),       //                                 .incoming_fifo_wrreq_signal
		.fee_2_rmap_outgoing_fifo_wrdata_flag_i (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal), //                                 .outgoing_fifo_wrdata_flag_signal
		.fee_2_rmap_outgoing_fifo_wrdata_data_i (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal), //                                 .outgoing_fifo_wrdata_data_signal
		.fee_2_rmap_outgoing_fifo_wrreq_i       (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal),       //                                 .outgoing_fifo_wrreq_signal
		.fee_3_rmap_echo_en_i                   (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_echo_en_signal),                   //   conduit_end_fee_3_rmap_echo_in.echo_en_signal
		.fee_3_rmap_echo_id_en_i                (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_echo_id_en_signal),                //                                 .echo_id_en_signal
		.fee_3_rmap_incoming_fifo_wrdata_flag_i (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal), //                                 .incoming_fifo_wrdata_flag_signal
		.fee_3_rmap_incoming_fifo_wrdata_data_i (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal), //                                 .incoming_fifo_wrdata_data_signal
		.fee_3_rmap_incoming_fifo_wrreq_i       (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal),       //                                 .incoming_fifo_wrreq_signal
		.fee_3_rmap_outgoing_fifo_wrdata_flag_i (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal), //                                 .outgoing_fifo_wrdata_flag_signal
		.fee_3_rmap_outgoing_fifo_wrdata_data_i (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal), //                                 .outgoing_fifo_wrdata_data_signal
		.fee_3_rmap_outgoing_fifo_wrreq_i       (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal),       //                                 .outgoing_fifo_wrreq_signal
		.fee_4_rmap_echo_en_i                   (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_echo_en_signal),                   //   conduit_end_fee_4_rmap_echo_in.echo_en_signal
		.fee_4_rmap_echo_id_en_i                (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_echo_id_en_signal),                //                                 .echo_id_en_signal
		.fee_4_rmap_incoming_fifo_wrdata_flag_i (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal), //                                 .incoming_fifo_wrdata_flag_signal
		.fee_4_rmap_incoming_fifo_wrdata_data_i (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal), //                                 .incoming_fifo_wrdata_data_signal
		.fee_4_rmap_incoming_fifo_wrreq_i       (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal),       //                                 .incoming_fifo_wrreq_signal
		.fee_4_rmap_outgoing_fifo_wrdata_flag_i (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal), //                                 .outgoing_fifo_wrdata_flag_signal
		.fee_4_rmap_outgoing_fifo_wrdata_data_i (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal), //                                 .outgoing_fifo_wrdata_data_signal
		.fee_4_rmap_outgoing_fifo_wrreq_i       (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal),       //                                 .outgoing_fifo_wrreq_signal
		.fee_5_rmap_echo_en_i                   (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_echo_en_signal),                   //   conduit_end_fee_5_rmap_echo_in.echo_en_signal
		.fee_5_rmap_echo_id_en_i                (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_echo_id_en_signal),                //                                 .echo_id_en_signal
		.fee_5_rmap_incoming_fifo_wrdata_flag_i (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_flag_signal), //                                 .incoming_fifo_wrdata_flag_signal
		.fee_5_rmap_incoming_fifo_wrdata_data_i (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_incoming_fifo_wrdata_data_signal), //                                 .incoming_fifo_wrdata_data_signal
		.fee_5_rmap_incoming_fifo_wrreq_i       (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_incoming_fifo_wrreq_signal),       //                                 .incoming_fifo_wrreq_signal
		.fee_5_rmap_outgoing_fifo_wrdata_flag_i (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_flag_signal), //                                 .outgoing_fifo_wrdata_flag_signal
		.fee_5_rmap_outgoing_fifo_wrdata_data_i (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrdata_data_signal), //                                 .outgoing_fifo_wrdata_data_signal
		.fee_5_rmap_outgoing_fifo_wrreq_i       (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_echo_out_outgoing_fifo_wrreq_signal),       //                                 .outgoing_fifo_wrreq_signal
		.spw_link_status_started_i              (spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_started_signal),     // conduit_end_spacewire_controller.spw_link_status_started_signal
		.spw_link_status_connecting_i           (spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_connecting_signal),  //                                 .spw_link_status_connecting_signal
		.spw_link_status_running_i              (spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_running_signal),     //                                 .spw_link_status_running_signal
		.spw_link_error_errdisc_i               (spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),      //                                 .spw_link_error_errdisc_signal
		.spw_link_error_errpar_i                (spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errpar_signal),       //                                 .spw_link_error_errpar_signal
		.spw_link_error_erresc_i                (spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_erresc_signal),       //                                 .spw_link_error_erresc_signal
		.spw_link_error_errcred_i               (spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errcred_signal),      //                                 .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_i             (spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),    //                                 .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_i             (spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),    //                                 .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_i             (spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),    //                                 .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_i           (spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),  //                                 .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_i           (spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),  //                                 .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_i            (spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),   //                                 .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_i            (spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),   //                                 .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_i             (spacewire_channel_h_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),    //                                 .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_i           (spacewire_channel_h_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal),  //                                 .spw_data_tx_status_txhalff_signal
		.spw_link_command_autostart_o           (rmap_echoing_0_conduit_end_spacewire_controller_spw_link_command_autostart_signal),    //                                 .spw_link_command_autostart_signal
		.spw_link_command_linkstart_o           (rmap_echoing_0_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),    //                                 .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_o             (rmap_echoing_0_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),      //                                 .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_o            (rmap_echoing_0_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),     //                                 .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_o              (rmap_echoing_0_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),       //                                 .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_o              (rmap_echoing_0_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),       //                                 .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_o              (rmap_echoing_0_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),       //                                 .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_o           (rmap_echoing_0_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),    //                                 .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_o          (rmap_echoing_0_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal),   //                                 .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_o           (rmap_echoing_0_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),    //                                 .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_o           (rmap_echoing_0_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal)     //                                 .spw_data_tx_command_txdata_signal
	);

	spwc_spacewire_channel_top spacewire_channel_a (
		.reset_i                       (rst_controller_010_reset_out_reset),                                                        //                    reset_sink.reset
		.clk_100_i                     (m2_ddr2_memory_afi_half_clk_clk),                                                           //             clock_sink_100mhz.clk
		.clk_200_i                     (m2_ddr2_memory_afi_clk_clk),                                                                //             clock_sink_200mhz.clk
		.spw_lvds_data_in_i            (spwc_a_lvds_spw_lvds_data_in_signal),                                                       //    conduit_end_spacewire_lvds.spw_lvds_data_in_signal
		.spw_lvds_data_out_o           (spwc_a_lvds_spw_lvds_data_out_signal),                                                      //                              .spw_lvds_data_out_signal
		.spw_lvds_strobe_out_o         (spwc_a_lvds_spw_lvds_strobe_out_signal),                                                    //                              .spw_lvds_strobe_out_signal
		.spw_lvds_strobe_in_i          (spwc_a_lvds_spw_lvds_strobe_in_signal),                                                     //                              .spw_lvds_strobe_in_signal
		.spw_rx_enable_i               (spwc_a_enable_spw_rx_enable_signal),                                                        //  conduit_end_spacewire_enable.spw_rx_enable_signal
		.spw_tx_enable_i               (spwc_a_enable_spw_tx_enable_signal),                                                        //                              .spw_tx_enable_signal
		.spw_red_status_led_o          (spwc_a_leds_spw_red_status_led_signal),                                                     //    conduit_end_spacewire_leds.spw_red_status_led_signal
		.spw_green_status_led_o        (spwc_a_leds_spw_green_status_led_signal),                                                   //                              .spw_green_status_led_signal
		.spw_link_command_autostart_i  (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_link_command_autostart_signal),  // conduit_end_spacewire_channel.spw_link_command_autostart_signal
		.spw_link_command_linkstart_i  (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),  //                              .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_i    (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),    //                              .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_i   (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),   //                              .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_i     (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),     //                              .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_i     (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),     //                              .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_i     (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),     //                              .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_i  (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),  //                              .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_i (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal), //                              .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_i  (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),  //                              .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_i  (comm_pedreiro_v1_01_1_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal),  //                              .spw_data_tx_command_txdata_signal
		.spw_link_status_started_o     (spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_started_signal),          //                              .spw_link_status_started_signal
		.spw_link_status_connecting_o  (spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_connecting_signal),       //                              .spw_link_status_connecting_signal
		.spw_link_status_running_o     (spacewire_channel_a_conduit_end_spacewire_channel_spw_link_status_running_signal),          //                              .spw_link_status_running_signal
		.spw_link_error_errdisc_o      (spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),           //                              .spw_link_error_errdisc_signal
		.spw_link_error_errpar_o       (spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errpar_signal),            //                              .spw_link_error_errpar_signal
		.spw_link_error_erresc_o       (spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_erresc_signal),            //                              .spw_link_error_erresc_signal
		.spw_link_error_errcred_o      (spacewire_channel_a_conduit_end_spacewire_channel_spw_link_error_errcred_signal),           //                              .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_o    (spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),         //                              .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_o    (spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),         //                              .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_o    (spacewire_channel_a_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),         //                              .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_o  (spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),       //                              .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_o  (spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),       //                              .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_o   (spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),        //                              .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_o   (spacewire_channel_a_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),        //                              .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_o    (spacewire_channel_a_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),         //                              .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_o  (spacewire_channel_a_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal)        //                              .spw_data_tx_status_txhalff_signal
	);

	spwc_spacewire_channel_top spacewire_channel_b (
		.reset_i                       (rst_controller_011_reset_out_reset),                                                        //                    reset_sink.reset
		.clk_100_i                     (m2_ddr2_memory_afi_half_clk_clk),                                                           //             clock_sink_100mhz.clk
		.clk_200_i                     (m2_ddr2_memory_afi_clk_clk),                                                                //             clock_sink_200mhz.clk
		.spw_lvds_data_in_i            (spwc_b_lvds_spw_lvds_data_in_signal),                                                       //    conduit_end_spacewire_lvds.spw_lvds_data_in_signal
		.spw_lvds_data_out_o           (spwc_b_lvds_spw_lvds_data_out_signal),                                                      //                              .spw_lvds_data_out_signal
		.spw_lvds_strobe_out_o         (spwc_b_lvds_spw_lvds_strobe_out_signal),                                                    //                              .spw_lvds_strobe_out_signal
		.spw_lvds_strobe_in_i          (spwc_b_lvds_spw_lvds_strobe_in_signal),                                                     //                              .spw_lvds_strobe_in_signal
		.spw_rx_enable_i               (spwc_b_enable_spw_rx_enable_signal),                                                        //  conduit_end_spacewire_enable.spw_rx_enable_signal
		.spw_tx_enable_i               (spwc_b_enable_spw_tx_enable_signal),                                                        //                              .spw_tx_enable_signal
		.spw_red_status_led_o          (spwc_b_leds_spw_red_status_led_signal),                                                     //    conduit_end_spacewire_leds.spw_red_status_led_signal
		.spw_green_status_led_o        (spwc_b_leds_spw_green_status_led_signal),                                                   //                              .spw_green_status_led_signal
		.spw_link_command_autostart_i  (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_link_command_autostart_signal),  // conduit_end_spacewire_channel.spw_link_command_autostart_signal
		.spw_link_command_linkstart_i  (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),  //                              .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_i    (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),    //                              .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_i   (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),   //                              .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_i     (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),     //                              .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_i     (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),     //                              .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_i     (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),     //                              .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_i  (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),  //                              .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_i (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal), //                              .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_i  (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),  //                              .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_i  (comm_pedreiro_v1_01_2_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal),  //                              .spw_data_tx_command_txdata_signal
		.spw_link_status_started_o     (spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_started_signal),          //                              .spw_link_status_started_signal
		.spw_link_status_connecting_o  (spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_connecting_signal),       //                              .spw_link_status_connecting_signal
		.spw_link_status_running_o     (spacewire_channel_b_conduit_end_spacewire_channel_spw_link_status_running_signal),          //                              .spw_link_status_running_signal
		.spw_link_error_errdisc_o      (spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),           //                              .spw_link_error_errdisc_signal
		.spw_link_error_errpar_o       (spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errpar_signal),            //                              .spw_link_error_errpar_signal
		.spw_link_error_erresc_o       (spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_erresc_signal),            //                              .spw_link_error_erresc_signal
		.spw_link_error_errcred_o      (spacewire_channel_b_conduit_end_spacewire_channel_spw_link_error_errcred_signal),           //                              .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_o    (spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),         //                              .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_o    (spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),         //                              .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_o    (spacewire_channel_b_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),         //                              .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_o  (spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),       //                              .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_o  (spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),       //                              .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_o   (spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),        //                              .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_o   (spacewire_channel_b_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),        //                              .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_o    (spacewire_channel_b_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),         //                              .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_o  (spacewire_channel_b_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal)        //                              .spw_data_tx_status_txhalff_signal
	);

	spwc_spacewire_channel_top spacewire_channel_c (
		.reset_i                       (rst_controller_012_reset_out_reset),                                                        //                    reset_sink.reset
		.clk_100_i                     (m2_ddr2_memory_afi_half_clk_clk),                                                           //             clock_sink_100mhz.clk
		.clk_200_i                     (m2_ddr2_memory_afi_clk_clk),                                                                //             clock_sink_200mhz.clk
		.spw_lvds_data_in_i            (spwc_c_lvds_spw_lvds_data_in_signal),                                                       //    conduit_end_spacewire_lvds.spw_lvds_data_in_signal
		.spw_lvds_data_out_o           (spwc_c_lvds_spw_lvds_data_out_signal),                                                      //                              .spw_lvds_data_out_signal
		.spw_lvds_strobe_out_o         (spwc_c_lvds_spw_lvds_strobe_out_signal),                                                    //                              .spw_lvds_strobe_out_signal
		.spw_lvds_strobe_in_i          (spwc_c_lvds_spw_lvds_strobe_in_signal),                                                     //                              .spw_lvds_strobe_in_signal
		.spw_rx_enable_i               (spwc_c_enable_spw_rx_enable_signal),                                                        //  conduit_end_spacewire_enable.spw_rx_enable_signal
		.spw_tx_enable_i               (spwc_c_enable_spw_tx_enable_signal),                                                        //                              .spw_tx_enable_signal
		.spw_red_status_led_o          (spwc_c_leds_spw_red_status_led_signal),                                                     //    conduit_end_spacewire_leds.spw_red_status_led_signal
		.spw_green_status_led_o        (spwc_c_leds_spw_green_status_led_signal),                                                   //                              .spw_green_status_led_signal
		.spw_link_command_autostart_i  (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_link_command_autostart_signal),  // conduit_end_spacewire_channel.spw_link_command_autostart_signal
		.spw_link_command_linkstart_i  (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),  //                              .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_i    (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),    //                              .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_i   (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),   //                              .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_i     (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),     //                              .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_i     (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),     //                              .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_i     (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),     //                              .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_i  (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),  //                              .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_i (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal), //                              .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_i  (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),  //                              .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_i  (comm_pedreiro_v1_01_3_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal),  //                              .spw_data_tx_command_txdata_signal
		.spw_link_status_started_o     (spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_started_signal),          //                              .spw_link_status_started_signal
		.spw_link_status_connecting_o  (spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_connecting_signal),       //                              .spw_link_status_connecting_signal
		.spw_link_status_running_o     (spacewire_channel_c_conduit_end_spacewire_channel_spw_link_status_running_signal),          //                              .spw_link_status_running_signal
		.spw_link_error_errdisc_o      (spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),           //                              .spw_link_error_errdisc_signal
		.spw_link_error_errpar_o       (spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errpar_signal),            //                              .spw_link_error_errpar_signal
		.spw_link_error_erresc_o       (spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_erresc_signal),            //                              .spw_link_error_erresc_signal
		.spw_link_error_errcred_o      (spacewire_channel_c_conduit_end_spacewire_channel_spw_link_error_errcred_signal),           //                              .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_o    (spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),         //                              .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_o    (spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),         //                              .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_o    (spacewire_channel_c_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),         //                              .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_o  (spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),       //                              .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_o  (spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),       //                              .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_o   (spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),        //                              .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_o   (spacewire_channel_c_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),        //                              .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_o    (spacewire_channel_c_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),         //                              .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_o  (spacewire_channel_c_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal)        //                              .spw_data_tx_status_txhalff_signal
	);

	spwc_spacewire_channel_top spacewire_channel_d (
		.reset_i                       (rst_controller_013_reset_out_reset),                                                        //                    reset_sink.reset
		.clk_100_i                     (m2_ddr2_memory_afi_half_clk_clk),                                                           //             clock_sink_100mhz.clk
		.clk_200_i                     (m2_ddr2_memory_afi_clk_clk),                                                                //             clock_sink_200mhz.clk
		.spw_lvds_data_in_i            (spwc_d_lvds_spw_lvds_data_in_signal),                                                       //    conduit_end_spacewire_lvds.spw_lvds_data_in_signal
		.spw_lvds_data_out_o           (spwc_d_lvds_spw_lvds_data_out_signal),                                                      //                              .spw_lvds_data_out_signal
		.spw_lvds_strobe_out_o         (spwc_d_lvds_spw_lvds_strobe_out_signal),                                                    //                              .spw_lvds_strobe_out_signal
		.spw_lvds_strobe_in_i          (spwc_d_lvds_spw_lvds_strobe_in_signal),                                                     //                              .spw_lvds_strobe_in_signal
		.spw_rx_enable_i               (spwc_d_enable_spw_rx_enable_signal),                                                        //  conduit_end_spacewire_enable.spw_rx_enable_signal
		.spw_tx_enable_i               (spwc_d_enable_spw_tx_enable_signal),                                                        //                              .spw_tx_enable_signal
		.spw_red_status_led_o          (spwc_d_leds_spw_red_status_led_signal),                                                     //    conduit_end_spacewire_leds.spw_red_status_led_signal
		.spw_green_status_led_o        (spwc_d_leds_spw_green_status_led_signal),                                                   //                              .spw_green_status_led_signal
		.spw_link_command_autostart_i  (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_link_command_autostart_signal),  // conduit_end_spacewire_channel.spw_link_command_autostart_signal
		.spw_link_command_linkstart_i  (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),  //                              .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_i    (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),    //                              .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_i   (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),   //                              .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_i     (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),     //                              .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_i     (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),     //                              .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_i     (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),     //                              .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_i  (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),  //                              .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_i (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal), //                              .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_i  (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),  //                              .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_i  (comm_pedreiro_v1_01_4_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal),  //                              .spw_data_tx_command_txdata_signal
		.spw_link_status_started_o     (spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_started_signal),          //                              .spw_link_status_started_signal
		.spw_link_status_connecting_o  (spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_connecting_signal),       //                              .spw_link_status_connecting_signal
		.spw_link_status_running_o     (spacewire_channel_d_conduit_end_spacewire_channel_spw_link_status_running_signal),          //                              .spw_link_status_running_signal
		.spw_link_error_errdisc_o      (spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),           //                              .spw_link_error_errdisc_signal
		.spw_link_error_errpar_o       (spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errpar_signal),            //                              .spw_link_error_errpar_signal
		.spw_link_error_erresc_o       (spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_erresc_signal),            //                              .spw_link_error_erresc_signal
		.spw_link_error_errcred_o      (spacewire_channel_d_conduit_end_spacewire_channel_spw_link_error_errcred_signal),           //                              .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_o    (spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),         //                              .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_o    (spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),         //                              .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_o    (spacewire_channel_d_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),         //                              .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_o  (spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),       //                              .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_o  (spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),       //                              .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_o   (spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),        //                              .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_o   (spacewire_channel_d_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),        //                              .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_o    (spacewire_channel_d_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),         //                              .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_o  (spacewire_channel_d_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal)        //                              .spw_data_tx_status_txhalff_signal
	);

	spwc_spacewire_channel_top spacewire_channel_e (
		.reset_i                       (rst_controller_014_reset_out_reset),                                                        //                    reset_sink.reset
		.clk_100_i                     (m2_ddr2_memory_afi_half_clk_clk),                                                           //             clock_sink_100mhz.clk
		.clk_200_i                     (m2_ddr2_memory_afi_clk_clk),                                                                //             clock_sink_200mhz.clk
		.spw_lvds_data_in_i            (spwc_e_lvds_spw_lvds_data_in_signal),                                                       //    conduit_end_spacewire_lvds.spw_lvds_data_in_signal
		.spw_lvds_data_out_o           (spwc_e_lvds_spw_lvds_data_out_signal),                                                      //                              .spw_lvds_data_out_signal
		.spw_lvds_strobe_out_o         (spwc_e_lvds_spw_lvds_strobe_out_signal),                                                    //                              .spw_lvds_strobe_out_signal
		.spw_lvds_strobe_in_i          (spwc_e_lvds_spw_lvds_strobe_in_signal),                                                     //                              .spw_lvds_strobe_in_signal
		.spw_rx_enable_i               (spwc_e_enable_spw_rx_enable_signal),                                                        //  conduit_end_spacewire_enable.spw_rx_enable_signal
		.spw_tx_enable_i               (spwc_e_enable_spw_tx_enable_signal),                                                        //                              .spw_tx_enable_signal
		.spw_red_status_led_o          (spwc_e_leds_spw_red_status_led_signal),                                                     //    conduit_end_spacewire_leds.spw_red_status_led_signal
		.spw_green_status_led_o        (spwc_e_leds_spw_green_status_led_signal),                                                   //                              .spw_green_status_led_signal
		.spw_link_command_autostart_i  (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_link_command_autostart_signal),  // conduit_end_spacewire_channel.spw_link_command_autostart_signal
		.spw_link_command_linkstart_i  (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),  //                              .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_i    (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),    //                              .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_i   (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),   //                              .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_i     (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),     //                              .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_i     (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),     //                              .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_i     (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),     //                              .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_i  (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),  //                              .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_i (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal), //                              .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_i  (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),  //                              .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_i  (comm_pedreiro_v1_01_5_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal),  //                              .spw_data_tx_command_txdata_signal
		.spw_link_status_started_o     (spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_started_signal),          //                              .spw_link_status_started_signal
		.spw_link_status_connecting_o  (spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_connecting_signal),       //                              .spw_link_status_connecting_signal
		.spw_link_status_running_o     (spacewire_channel_e_conduit_end_spacewire_channel_spw_link_status_running_signal),          //                              .spw_link_status_running_signal
		.spw_link_error_errdisc_o      (spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),           //                              .spw_link_error_errdisc_signal
		.spw_link_error_errpar_o       (spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errpar_signal),            //                              .spw_link_error_errpar_signal
		.spw_link_error_erresc_o       (spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_erresc_signal),            //                              .spw_link_error_erresc_signal
		.spw_link_error_errcred_o      (spacewire_channel_e_conduit_end_spacewire_channel_spw_link_error_errcred_signal),           //                              .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_o    (spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),         //                              .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_o    (spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),         //                              .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_o    (spacewire_channel_e_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),         //                              .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_o  (spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),       //                              .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_o  (spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),       //                              .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_o   (spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),        //                              .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_o   (spacewire_channel_e_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),        //                              .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_o    (spacewire_channel_e_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),         //                              .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_o  (spacewire_channel_e_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal)        //                              .spw_data_tx_status_txhalff_signal
	);

	spwc_spacewire_channel_top spacewire_channel_f (
		.reset_i                       (rst_controller_015_reset_out_reset),                                                        //                    reset_sink.reset
		.clk_100_i                     (m2_ddr2_memory_afi_half_clk_clk),                                                           //             clock_sink_100mhz.clk
		.clk_200_i                     (m2_ddr2_memory_afi_clk_clk),                                                                //             clock_sink_200mhz.clk
		.spw_lvds_data_in_i            (spwc_f_lvds_spw_lvds_data_in_signal),                                                       //    conduit_end_spacewire_lvds.spw_lvds_data_in_signal
		.spw_lvds_data_out_o           (spwc_f_lvds_spw_lvds_data_out_signal),                                                      //                              .spw_lvds_data_out_signal
		.spw_lvds_strobe_out_o         (spwc_f_lvds_spw_lvds_strobe_out_signal),                                                    //                              .spw_lvds_strobe_out_signal
		.spw_lvds_strobe_in_i          (spwc_f_lvds_spw_lvds_strobe_in_signal),                                                     //                              .spw_lvds_strobe_in_signal
		.spw_rx_enable_i               (spwc_f_enable_spw_rx_enable_signal),                                                        //  conduit_end_spacewire_enable.spw_rx_enable_signal
		.spw_tx_enable_i               (spwc_f_enable_spw_tx_enable_signal),                                                        //                              .spw_tx_enable_signal
		.spw_red_status_led_o          (spwc_f_leds_spw_red_status_led_signal),                                                     //    conduit_end_spacewire_leds.spw_red_status_led_signal
		.spw_green_status_led_o        (spwc_f_leds_spw_green_status_led_signal),                                                   //                              .spw_green_status_led_signal
		.spw_link_command_autostart_i  (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_link_command_autostart_signal),  // conduit_end_spacewire_channel.spw_link_command_autostart_signal
		.spw_link_command_linkstart_i  (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),  //                              .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_i    (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),    //                              .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_i   (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),   //                              .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_i     (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),     //                              .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_i     (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),     //                              .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_i     (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),     //                              .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_i  (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),  //                              .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_i (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal), //                              .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_i  (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),  //                              .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_i  (comm_pedreiro_v1_01_6_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal),  //                              .spw_data_tx_command_txdata_signal
		.spw_link_status_started_o     (spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_started_signal),          //                              .spw_link_status_started_signal
		.spw_link_status_connecting_o  (spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_connecting_signal),       //                              .spw_link_status_connecting_signal
		.spw_link_status_running_o     (spacewire_channel_f_conduit_end_spacewire_channel_spw_link_status_running_signal),          //                              .spw_link_status_running_signal
		.spw_link_error_errdisc_o      (spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),           //                              .spw_link_error_errdisc_signal
		.spw_link_error_errpar_o       (spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errpar_signal),            //                              .spw_link_error_errpar_signal
		.spw_link_error_erresc_o       (spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_erresc_signal),            //                              .spw_link_error_erresc_signal
		.spw_link_error_errcred_o      (spacewire_channel_f_conduit_end_spacewire_channel_spw_link_error_errcred_signal),           //                              .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_o    (spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),         //                              .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_o    (spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),         //                              .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_o    (spacewire_channel_f_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),         //                              .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_o  (spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),       //                              .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_o  (spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),       //                              .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_o   (spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),        //                              .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_o   (spacewire_channel_f_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),        //                              .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_o    (spacewire_channel_f_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),         //                              .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_o  (spacewire_channel_f_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal)        //                              .spw_data_tx_status_txhalff_signal
	);

	spwc_spacewire_channel_top spacewire_channel_g (
		.reset_i                       (rst_controller_016_reset_out_reset),                                                      //                    reset_sink.reset
		.clk_100_i                     (m2_ddr2_memory_afi_half_clk_clk),                                                         //             clock_sink_100mhz.clk
		.clk_200_i                     (m2_ddr2_memory_afi_clk_clk),                                                              //             clock_sink_200mhz.clk
		.spw_lvds_data_in_i            (spwc_g_lvds_spw_lvds_data_in_signal),                                                     //    conduit_end_spacewire_lvds.spw_lvds_data_in_signal
		.spw_lvds_data_out_o           (spwc_g_lvds_spw_lvds_data_out_signal),                                                    //                              .spw_lvds_data_out_signal
		.spw_lvds_strobe_out_o         (spwc_g_lvds_spw_lvds_strobe_out_signal),                                                  //                              .spw_lvds_strobe_out_signal
		.spw_lvds_strobe_in_i          (spwc_g_lvds_spw_lvds_strobe_in_signal),                                                   //                              .spw_lvds_strobe_in_signal
		.spw_rx_enable_i               (spwc_g_enable_spw_rx_enable_signal),                                                      //  conduit_end_spacewire_enable.spw_rx_enable_signal
		.spw_tx_enable_i               (spwc_g_enable_spw_tx_enable_signal),                                                      //                              .spw_tx_enable_signal
		.spw_red_status_led_o          (spwc_g_leds_spw_red_status_led_signal),                                                   //    conduit_end_spacewire_leds.spw_red_status_led_signal
		.spw_green_status_led_o        (spwc_g_leds_spw_green_status_led_signal),                                                 //                              .spw_green_status_led_signal
		.spw_link_command_autostart_i  (spacewire_glutton_0_conduit_end_spacewire_controller_spw_link_command_autostart_signal),  // conduit_end_spacewire_channel.spw_link_command_autostart_signal
		.spw_link_command_linkstart_i  (spacewire_glutton_0_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),  //                              .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_i    (spacewire_glutton_0_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),    //                              .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_i   (spacewire_glutton_0_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),   //                              .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_i     (spacewire_glutton_0_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),     //                              .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_i     (spacewire_glutton_0_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),     //                              .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_i     (spacewire_glutton_0_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),     //                              .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_i  (spacewire_glutton_0_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),  //                              .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_i (spacewire_glutton_0_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal), //                              .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_i  (spacewire_glutton_0_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),  //                              .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_i  (spacewire_glutton_0_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal),  //                              .spw_data_tx_command_txdata_signal
		.spw_link_status_started_o     (spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_started_signal),        //                              .spw_link_status_started_signal
		.spw_link_status_connecting_o  (spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_connecting_signal),     //                              .spw_link_status_connecting_signal
		.spw_link_status_running_o     (spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_running_signal),        //                              .spw_link_status_running_signal
		.spw_link_error_errdisc_o      (spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),         //                              .spw_link_error_errdisc_signal
		.spw_link_error_errpar_o       (spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errpar_signal),          //                              .spw_link_error_errpar_signal
		.spw_link_error_erresc_o       (spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_erresc_signal),          //                              .spw_link_error_erresc_signal
		.spw_link_error_errcred_o      (spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errcred_signal),         //                              .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_o    (spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),       //                              .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_o    (spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),       //                              .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_o    (spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),       //                              .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_o  (spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),     //                              .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_o  (spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),     //                              .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_o   (spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),      //                              .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_o   (spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),      //                              .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_o    (spacewire_channel_g_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),       //                              .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_o  (spacewire_channel_g_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal)      //                              .spw_data_tx_status_txhalff_signal
	);

	spwc_spacewire_channel_top spacewire_channel_h (
		.reset_i                       (rst_controller_017_reset_out_reset),                                                  //                    reset_sink.reset
		.clk_100_i                     (m2_ddr2_memory_afi_half_clk_clk),                                                     //             clock_sink_100mhz.clk
		.clk_200_i                     (m2_ddr2_memory_afi_clk_clk),                                                          //             clock_sink_200mhz.clk
		.spw_lvds_data_in_i            (spwc_h_lvds_spw_lvds_data_in_signal),                                                 //    conduit_end_spacewire_lvds.spw_lvds_data_in_signal
		.spw_lvds_data_out_o           (spwc_h_lvds_spw_lvds_data_out_signal),                                                //                              .spw_lvds_data_out_signal
		.spw_lvds_strobe_out_o         (spwc_h_lvds_spw_lvds_strobe_out_signal),                                              //                              .spw_lvds_strobe_out_signal
		.spw_lvds_strobe_in_i          (spwc_h_lvds_spw_lvds_strobe_in_signal),                                               //                              .spw_lvds_strobe_in_signal
		.spw_rx_enable_i               (spwc_h_enable_spw_rx_enable_signal),                                                  //  conduit_end_spacewire_enable.spw_rx_enable_signal
		.spw_tx_enable_i               (spwc_h_enable_spw_tx_enable_signal),                                                  //                              .spw_tx_enable_signal
		.spw_red_status_led_o          (spwc_h_leds_spw_red_status_led_signal),                                               //    conduit_end_spacewire_leds.spw_red_status_led_signal
		.spw_green_status_led_o        (spwc_h_leds_spw_green_status_led_signal),                                             //                              .spw_green_status_led_signal
		.spw_link_command_autostart_i  (rmap_echoing_0_conduit_end_spacewire_controller_spw_link_command_autostart_signal),   // conduit_end_spacewire_channel.spw_link_command_autostart_signal
		.spw_link_command_linkstart_i  (rmap_echoing_0_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),   //                              .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_i    (rmap_echoing_0_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),     //                              .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_i   (rmap_echoing_0_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),    //                              .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_i     (rmap_echoing_0_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),      //                              .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_i     (rmap_echoing_0_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),      //                              .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_i     (rmap_echoing_0_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),      //                              .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_i  (rmap_echoing_0_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),   //                              .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_i (rmap_echoing_0_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal),  //                              .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_i  (rmap_echoing_0_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),   //                              .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_i  (rmap_echoing_0_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal),   //                              .spw_data_tx_command_txdata_signal
		.spw_link_status_started_o     (spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_started_signal),    //                              .spw_link_status_started_signal
		.spw_link_status_connecting_o  (spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_connecting_signal), //                              .spw_link_status_connecting_signal
		.spw_link_status_running_o     (spacewire_channel_h_conduit_end_spacewire_channel_spw_link_status_running_signal),    //                              .spw_link_status_running_signal
		.spw_link_error_errdisc_o      (spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),     //                              .spw_link_error_errdisc_signal
		.spw_link_error_errpar_o       (spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errpar_signal),      //                              .spw_link_error_errpar_signal
		.spw_link_error_erresc_o       (spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_erresc_signal),      //                              .spw_link_error_erresc_signal
		.spw_link_error_errcred_o      (spacewire_channel_h_conduit_end_spacewire_channel_spw_link_error_errcred_signal),     //                              .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_o    (spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),   //                              .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_o    (spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),   //                              .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_o    (spacewire_channel_h_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),   //                              .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_o  (spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal), //                              .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_o  (spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal), //                              .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_o   (spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),  //                              .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_o   (spacewire_channel_h_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),  //                              .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_o    (spacewire_channel_h_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),   //                              .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_o  (spacewire_channel_h_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal)  //                              .spw_data_tx_status_txhalff_signal
	);

	spwg_spw_glutton_top spacewire_glutton_0 (
		.reset_i                       (rst_controller_018_reset_out_reset),                                                      //                       reset_sink.reset
		.clk_100_i                     (m2_ddr2_memory_afi_half_clk_clk),                                                         //                clock_sink_100mhz.clk
		.spw_link_status_started_i     (spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_started_signal),        // conduit_end_spacewire_controller.spw_link_status_started_signal
		.spw_link_status_connecting_i  (spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_connecting_signal),     //                                 .spw_link_status_connecting_signal
		.spw_link_status_running_i     (spacewire_channel_g_conduit_end_spacewire_channel_spw_link_status_running_signal),        //                                 .spw_link_status_running_signal
		.spw_link_error_errdisc_i      (spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errdisc_signal),         //                                 .spw_link_error_errdisc_signal
		.spw_link_error_errpar_i       (spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errpar_signal),          //                                 .spw_link_error_errpar_signal
		.spw_link_error_erresc_i       (spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_erresc_signal),          //                                 .spw_link_error_erresc_signal
		.spw_link_error_errcred_i      (spacewire_channel_g_conduit_end_spacewire_channel_spw_link_error_errcred_signal),         //                                 .spw_link_error_errcred_signal
		.spw_timecode_rx_tick_out_i    (spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_tick_out_signal),       //                                 .spw_timecode_rx_tick_out_signal
		.spw_timecode_rx_ctrl_out_i    (spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_ctrl_out_signal),       //                                 .spw_timecode_rx_ctrl_out_signal
		.spw_timecode_rx_time_out_i    (spacewire_channel_g_conduit_end_spacewire_channel_spw_timecode_rx_time_out_signal),       //                                 .spw_timecode_rx_time_out_signal
		.spw_data_rx_status_rxvalid_i  (spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxvalid_signal),     //                                 .spw_data_rx_status_rxvalid_signal
		.spw_data_rx_status_rxhalff_i  (spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxhalff_signal),     //                                 .spw_data_rx_status_rxhalff_signal
		.spw_data_rx_status_rxflag_i   (spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxflag_signal),      //                                 .spw_data_rx_status_rxflag_signal
		.spw_data_rx_status_rxdata_i   (spacewire_channel_g_conduit_end_spacewire_channel_spw_data_rx_status_rxdata_signal),      //                                 .spw_data_rx_status_rxdata_signal
		.spw_data_tx_status_txrdy_i    (spacewire_channel_g_conduit_end_spacewire_channel_spw_data_tx_status_txrdy_signal),       //                                 .spw_data_tx_status_txrdy_signal
		.spw_data_tx_status_txhalff_i  (spacewire_channel_g_conduit_end_spacewire_channel_spw_data_tx_status_txhalff_signal),     //                                 .spw_data_tx_status_txhalff_signal
		.spw_link_command_autostart_o  (spacewire_glutton_0_conduit_end_spacewire_controller_spw_link_command_autostart_signal),  //                                 .spw_link_command_autostart_signal
		.spw_link_command_linkstart_o  (spacewire_glutton_0_conduit_end_spacewire_controller_spw_link_command_linkstart_signal),  //                                 .spw_link_command_linkstart_signal
		.spw_link_command_linkdis_o    (spacewire_glutton_0_conduit_end_spacewire_controller_spw_link_command_linkdis_signal),    //                                 .spw_link_command_linkdis_signal
		.spw_link_command_txdivcnt_o   (spacewire_glutton_0_conduit_end_spacewire_controller_spw_link_command_txdivcnt_signal),   //                                 .spw_link_command_txdivcnt_signal
		.spw_timecode_tx_tick_in_o     (spacewire_glutton_0_conduit_end_spacewire_controller_spw_timecode_tx_tick_in_signal),     //                                 .spw_timecode_tx_tick_in_signal
		.spw_timecode_tx_ctrl_in_o     (spacewire_glutton_0_conduit_end_spacewire_controller_spw_timecode_tx_ctrl_in_signal),     //                                 .spw_timecode_tx_ctrl_in_signal
		.spw_timecode_tx_time_in_o     (spacewire_glutton_0_conduit_end_spacewire_controller_spw_timecode_tx_time_in_signal),     //                                 .spw_timecode_tx_time_in_signal
		.spw_data_rx_command_rxread_o  (spacewire_glutton_0_conduit_end_spacewire_controller_spw_data_rx_command_rxread_signal),  //                                 .spw_data_rx_command_rxread_signal
		.spw_data_tx_command_txwrite_o (spacewire_glutton_0_conduit_end_spacewire_controller_spw_data_tx_command_txwrite_signal), //                                 .spw_data_tx_command_txwrite_signal
		.spw_data_tx_command_txflag_o  (spacewire_glutton_0_conduit_end_spacewire_controller_spw_data_tx_command_txflag_signal),  //                                 .spw_data_tx_command_txflag_signal
		.spw_data_tx_command_txdata_o  (spacewire_glutton_0_conduit_end_spacewire_controller_spw_data_tx_command_txdata_signal)   //                                 .spw_data_tx_command_txdata_signal
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (12),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) clock_bridge_afi_50 (
		.m0_clk           (clk50_clk),                                              //   m0_clk.clk
		.m0_reset         (rst_controller_019_reset_out_reset),                     // m0_reset.reset
		.s0_clk           (m2_ddr2_memory_afi_half_clk_clk),                        //   s0_clk.clk
		.s0_reset         (rst_controller_008_reset_out_reset),                     // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_1_clock_bridge_afi_50_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_1_clock_bridge_afi_50_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_1_clock_bridge_afi_50_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_1_clock_bridge_afi_50_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_1_clock_bridge_afi_50_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_1_clock_bridge_afi_50_s0_address),       //         .address
		.s0_write         (mm_interconnect_1_clock_bridge_afi_50_s0_write),         //         .write
		.s0_read          (mm_interconnect_1_clock_bridge_afi_50_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_1_clock_bridge_afi_50_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_1_clock_bridge_afi_50_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_bridge_afi_50_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_bridge_afi_50_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_bridge_afi_50_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_bridge_afi_50_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_bridge_afi_50_m0_writedata),                       //         .writedata
		.m0_address       (clock_bridge_afi_50_m0_address),                         //         .address
		.m0_write         (clock_bridge_afi_50_m0_write),                           //         .write
		.m0_read          (clock_bridge_afi_50_m0_read),                            //         .read
		.m0_byteenable    (clock_bridge_afi_50_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_bridge_afi_50_m0_debugaccess)                      //         .debugaccess
	);

	MebX_Qsys_Project_csense_adc_fo csense_adc_fo (
		.clk        (clk50_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_2_csense_adc_fo_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_csense_adc_fo_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_csense_adc_fo_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_csense_adc_fo_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_csense_adc_fo_s1_readdata),   //                    .readdata
		.out_port   (csense_adc_fo_export)                           // external_connection.export
	);

	MebX_Qsys_Project_csense_cs_n csense_cs_n (
		.clk        (clk50_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_2_csense_cs_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_csense_cs_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_csense_cs_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_csense_cs_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_csense_cs_n_s1_readdata),   //                    .readdata
		.out_port   (csense_cs_n_export)                           // external_connection.export
	);

	MebX_Qsys_Project_csense_adc_fo csense_sck (
		.clk        (clk50_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_2_csense_sck_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_csense_sck_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_csense_sck_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_csense_sck_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_csense_sck_s1_readdata),   //                    .readdata
		.out_port   (csense_sck_export)                           // external_connection.export
	);

	MebX_Qsys_Project_csense_adc_fo csense_sdi (
		.clk        (clk50_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_2_csense_sdi_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_csense_sdi_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_csense_sdi_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_csense_sdi_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_csense_sdi_s1_readdata),   //                    .readdata
		.out_port   (csense_sdi_export)                           // external_connection.export
	);

	MebX_Qsys_Project_csense_sdo csense_sdo (
		.clk      (clk50_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_019_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_2_csense_sdo_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_csense_sdo_s1_readdata), //                    .readdata
		.in_port  (csense_sdo_export)                         // external_connection.export
	);

	altera_address_span_extender #(
		.DATA_WIDTH           (32),
		.BYTEENABLE_WIDTH     (4),
		.MASTER_ADDRESS_WIDTH (32),
		.SLAVE_ADDRESS_WIDTH  (29),
		.SLAVE_ADDRESS_SHIFT  (2),
		.BURSTCOUNT_WIDTH     (8),
		.CNTL_ADDRESS_WIDTH   (1),
		.SUB_WINDOW_COUNT     (1),
		.MASTER_ADDRESS_DEF   (64'b0000000000000000000000000000000000000000000000000000000000000000)
	) ddr2_address_span_extender (
		.clk                  (m2_ddr2_memory_afi_half_clk_clk),                                           //           clock.clk
		.reset                (rst_controller_008_reset_out_reset),                                        //           reset.reset
		.avs_s0_address       (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_address),       //  windowed_slave.address
		.avs_s0_read          (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_read),          //                .read
		.avs_s0_readdata      (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdata),      //                .readdata
		.avs_s0_write         (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_write),         //                .write
		.avs_s0_writedata     (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_writedata),     //                .writedata
		.avs_s0_readdatavalid (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdatavalid), //                .readdatavalid
		.avs_s0_waitrequest   (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_waitrequest),   //                .waitrequest
		.avs_s0_byteenable    (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_byteenable),    //                .byteenable
		.avs_s0_burstcount    (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_burstcount),    //                .burstcount
		.avm_m0_address       (ddr2_address_span_extender_expanded_master_address),                        // expanded_master.address
		.avm_m0_read          (ddr2_address_span_extender_expanded_master_read),                           //                .read
		.avm_m0_waitrequest   (ddr2_address_span_extender_expanded_master_waitrequest),                    //                .waitrequest
		.avm_m0_readdata      (ddr2_address_span_extender_expanded_master_readdata),                       //                .readdata
		.avm_m0_write         (ddr2_address_span_extender_expanded_master_write),                          //                .write
		.avm_m0_writedata     (ddr2_address_span_extender_expanded_master_writedata),                      //                .writedata
		.avm_m0_readdatavalid (ddr2_address_span_extender_expanded_master_readdatavalid),                  //                .readdatavalid
		.avm_m0_byteenable    (ddr2_address_span_extender_expanded_master_byteenable),                     //                .byteenable
		.avm_m0_burstcount    (ddr2_address_span_extender_expanded_master_burstcount),                     //                .burstcount
		.avs_cntl_read        (mm_interconnect_1_ddr2_address_span_extender_cntl_read),                    //            cntl.read
		.avs_cntl_readdata    (mm_interconnect_1_ddr2_address_span_extender_cntl_readdata),                //                .readdata
		.avs_cntl_write       (mm_interconnect_1_ddr2_address_span_extender_cntl_write),                   //                .write
		.avs_cntl_writedata   (mm_interconnect_1_ddr2_address_span_extender_cntl_writedata),               //                .writedata
		.avs_cntl_byteenable  (mm_interconnect_1_ddr2_address_span_extender_cntl_byteenable),              //                .byteenable
		.avs_cntl_address     (1'b0)                                                                       //     (terminated)
	);

	MebX_Qsys_Project_ext_flash #(
		.TCM_ADDRESS_W                  (26),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (100),
		.TCM_WRITE_WAIT                 (100),
		.TCM_SETUP_WAIT                 (25),
		.TCM_DATA_HOLD                  (20),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) ext_flash (
		.clk_clk              (m2_ddr2_memory_afi_half_clk_clk),               //   clk.clk
		.reset_reset          (rst_controller_020_reset_out_reset),            // reset.reset
		.uas_address          (mm_interconnect_1_ext_flash_uas_address),       //   uas.address
		.uas_burstcount       (mm_interconnect_1_ext_flash_uas_burstcount),    //      .burstcount
		.uas_read             (mm_interconnect_1_ext_flash_uas_read),          //      .read
		.uas_write            (mm_interconnect_1_ext_flash_uas_write),         //      .write
		.uas_waitrequest      (mm_interconnect_1_ext_flash_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (mm_interconnect_1_ext_flash_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable       (mm_interconnect_1_ext_flash_uas_byteenable),    //      .byteenable
		.uas_readdata         (mm_interconnect_1_ext_flash_uas_readdata),      //      .readdata
		.uas_writedata        (mm_interconnect_1_ext_flash_uas_writedata),     //      .writedata
		.uas_lock             (mm_interconnect_1_ext_flash_uas_lock),          //      .lock
		.uas_debugaccess      (mm_interconnect_1_ext_flash_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (ext_flash_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_read_n_out       (ext_flash_tcm_read_n_out),                      //      .read_n_out
		.tcm_chipselect_n_out (ext_flash_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_request          (ext_flash_tcm_request),                         //      .request
		.tcm_grant            (ext_flash_tcm_grant),                           //      .grant
		.tcm_address_out      (ext_flash_tcm_address_out),                     //      .address_out
		.tcm_data_out         (ext_flash_tcm_data_out),                        //      .data_out
		.tcm_data_outen       (ext_flash_tcm_data_outen),                      //      .data_outen
		.tcm_data_in          (ext_flash_tcm_data_in)                          //      .data_in
	);

	MebX_Qsys_Project_jtag_uart_0 jtag_uart_0 (
		.clk            (m2_ddr2_memory_afi_half_clk_clk),                             //               clk.clk
		.rst_n          (~rst_controller_008_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver8_irq)                                     //               irq.irq
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (256),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (31),
		.BURSTCOUNT_WIDTH    (3),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (8),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) m1_clock_bridge (
		.m0_clk           (m1_ddr2_memory_afi_half_clk_clk),                    //   m0_clk.clk
		.m0_reset         (rst_controller_021_reset_out_reset),                 // m0_reset.reset
		.s0_clk           (m2_ddr2_memory_afi_half_clk_clk),                    //   s0_clk.clk
		.s0_reset         (rst_controller_008_reset_out_reset),                 // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_m1_clock_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_m1_clock_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_m1_clock_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_m1_clock_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_m1_clock_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_m1_clock_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_m1_clock_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_m1_clock_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_m1_clock_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_m1_clock_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (m1_clock_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (m1_clock_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (m1_clock_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (m1_clock_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (m1_clock_bridge_m0_writedata),                       //         .writedata
		.m0_address       (m1_clock_bridge_m0_address),                         //         .address
		.m0_write         (m1_clock_bridge_m0_write),                           //         .write
		.m0_read          (m1_clock_bridge_m0_read),                            //         .read
		.m0_byteenable    (m1_clock_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (m1_clock_bridge_m0_debugaccess)                      //         .debugaccess
	);

	MebX_Qsys_Project_csense_adc_fo m1_ddr2_i2c_scl (
		.clk        (clk50_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_2_m1_ddr2_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_m1_ddr2_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_m1_ddr2_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_m1_ddr2_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_m1_ddr2_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (m1_ddr2_i2c_scl_export)                           // external_connection.export
	);

	MebX_Qsys_Project_m1_ddr2_i2c_sda m1_ddr2_i2c_sda (
		.clk        (clk50_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_2_m1_ddr2_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_m1_ddr2_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_m1_ddr2_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_m1_ddr2_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_m1_ddr2_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (m1_ddr2_i2c_sda_export)                           // external_connection.export
	);

	MebX_Qsys_Project_m1_ddr2_memory m1_ddr2_memory (
		.pll_ref_clk        (m1_ddr2_memory_pll_ref_clk_clk),                          //      pll_ref_clk.clk
		.global_reset_n     (rst_reset_n),                                             //     global_reset.reset_n
		.soft_reset_n       (rst_reset_n),                                             //       soft_reset.reset_n
		.afi_clk            (m1_ddr2_memory_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk       (m1_ddr2_memory_afi_half_clk_clk),                         //     afi_half_clk.clk
		.afi_reset_n        (),                                                        //        afi_reset.reset_n
		.afi_reset_export_n (),                                                        // afi_reset_export.reset_n
		.mem_a              (m1_ddr2_memory_mem_a),                                    //           memory.mem_a
		.mem_ba             (m1_ddr2_memory_mem_ba),                                   //                 .mem_ba
		.mem_ck             (m1_ddr2_memory_mem_ck),                                   //                 .mem_ck
		.mem_ck_n           (m1_ddr2_memory_mem_ck_n),                                 //                 .mem_ck_n
		.mem_cke            (m1_ddr2_memory_mem_cke),                                  //                 .mem_cke
		.mem_cs_n           (m1_ddr2_memory_mem_cs_n),                                 //                 .mem_cs_n
		.mem_dm             (m1_ddr2_memory_mem_dm),                                   //                 .mem_dm
		.mem_ras_n          (m1_ddr2_memory_mem_ras_n),                                //                 .mem_ras_n
		.mem_cas_n          (m1_ddr2_memory_mem_cas_n),                                //                 .mem_cas_n
		.mem_we_n           (m1_ddr2_memory_mem_we_n),                                 //                 .mem_we_n
		.mem_dq             (m1_ddr2_memory_mem_dq),                                   //                 .mem_dq
		.mem_dqs            (m1_ddr2_memory_mem_dqs),                                  //                 .mem_dqs
		.mem_dqs_n          (m1_ddr2_memory_mem_dqs_n),                                //                 .mem_dqs_n
		.mem_odt            (m1_ddr2_memory_mem_odt),                                  //                 .mem_odt
		.avl_ready          (mm_interconnect_3_m1_ddr2_memory_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin     (mm_interconnect_3_m1_ddr2_memory_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr           (mm_interconnect_3_m1_ddr2_memory_avl_address),            //                 .address
		.avl_rdata_valid    (mm_interconnect_3_m1_ddr2_memory_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata          (mm_interconnect_3_m1_ddr2_memory_avl_readdata),           //                 .readdata
		.avl_wdata          (mm_interconnect_3_m1_ddr2_memory_avl_writedata),          //                 .writedata
		.avl_be             (mm_interconnect_3_m1_ddr2_memory_avl_byteenable),         //                 .byteenable
		.avl_read_req       (mm_interconnect_3_m1_ddr2_memory_avl_read),               //                 .read
		.avl_write_req      (mm_interconnect_3_m1_ddr2_memory_avl_write),              //                 .write
		.avl_size           (mm_interconnect_3_m1_ddr2_memory_avl_burstcount),         //                 .burstcount
		.local_init_done    (m1_ddr2_memory_status_local_init_done),                   //           status.local_init_done
		.local_cal_success  (m1_ddr2_memory_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail     (m1_ddr2_memory_status_local_cal_fail),                    //                 .local_cal_fail
		.oct_rdn            (m1_ddr2_oct_rdn),                                         //              oct.rdn
		.oct_rup            (m1_ddr2_oct_rup)                                          //                 .rup
	);

	MebX_Qsys_Project_csense_adc_fo m2_ddr2_i2c_scl (
		.clk        (clk50_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_2_m2_ddr2_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_m2_ddr2_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_m2_ddr2_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_m2_ddr2_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_m2_ddr2_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (m2_ddr2_i2c_scl_export)                           // external_connection.export
	);

	MebX_Qsys_Project_m1_ddr2_i2c_sda m2_ddr2_i2c_sda (
		.clk        (clk50_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_2_m2_ddr2_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_m2_ddr2_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_m2_ddr2_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_m2_ddr2_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_m2_ddr2_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (m2_ddr2_i2c_sda_export)                           // external_connection.export
	);

	MebX_Qsys_Project_m2_ddr2_memory m2_ddr2_memory (
		.pll_ref_clk               (clk50_clk),                                               //      pll_ref_clk.clk
		.global_reset_n            (rst_reset_n),                                             //     global_reset.reset_n
		.soft_reset_n              (rst_reset_n),                                             //       soft_reset.reset_n
		.afi_clk                   (m2_ddr2_memory_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk              (m2_ddr2_memory_afi_half_clk_clk),                         //     afi_half_clk.clk
		.afi_reset_n               (),                                                        //        afi_reset.reset_n
		.afi_reset_export_n        (),                                                        // afi_reset_export.reset_n
		.mem_a                     (m2_ddr2_memory_mem_a),                                    //           memory.mem_a
		.mem_ba                    (m2_ddr2_memory_mem_ba),                                   //                 .mem_ba
		.mem_ck                    (m2_ddr2_memory_mem_ck),                                   //                 .mem_ck
		.mem_ck_n                  (m2_ddr2_memory_mem_ck_n),                                 //                 .mem_ck_n
		.mem_cke                   (m2_ddr2_memory_mem_cke),                                  //                 .mem_cke
		.mem_cs_n                  (m2_ddr2_memory_mem_cs_n),                                 //                 .mem_cs_n
		.mem_dm                    (m2_ddr2_memory_mem_dm),                                   //                 .mem_dm
		.mem_ras_n                 (m2_ddr2_memory_mem_ras_n),                                //                 .mem_ras_n
		.mem_cas_n                 (m2_ddr2_memory_mem_cas_n),                                //                 .mem_cas_n
		.mem_we_n                  (m2_ddr2_memory_mem_we_n),                                 //                 .mem_we_n
		.mem_dq                    (m2_ddr2_memory_mem_dq),                                   //                 .mem_dq
		.mem_dqs                   (m2_ddr2_memory_mem_dqs),                                  //                 .mem_dqs
		.mem_dqs_n                 (m2_ddr2_memory_mem_dqs_n),                                //                 .mem_dqs_n
		.mem_odt                   (m2_ddr2_memory_mem_odt),                                  //                 .mem_odt
		.avl_ready                 (mm_interconnect_0_m2_ddr2_memory_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin            (mm_interconnect_0_m2_ddr2_memory_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (mm_interconnect_0_m2_ddr2_memory_avl_address),            //                 .address
		.avl_rdata_valid           (mm_interconnect_0_m2_ddr2_memory_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (mm_interconnect_0_m2_ddr2_memory_avl_readdata),           //                 .readdata
		.avl_wdata                 (mm_interconnect_0_m2_ddr2_memory_avl_writedata),          //                 .writedata
		.avl_be                    (mm_interconnect_0_m2_ddr2_memory_avl_byteenable),         //                 .byteenable
		.avl_read_req              (mm_interconnect_0_m2_ddr2_memory_avl_read),               //                 .read
		.avl_write_req             (mm_interconnect_0_m2_ddr2_memory_avl_write),              //                 .write
		.avl_size                  (mm_interconnect_0_m2_ddr2_memory_avl_burstcount),         //                 .burstcount
		.local_init_done           (m2_ddr2_memory_status_local_init_done),                   //           status.local_init_done
		.local_cal_success         (m2_ddr2_memory_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail            (m2_ddr2_memory_status_local_cal_fail),                    //                 .local_cal_fail
		.oct_rdn                   (m2_ddr2_oct_rdn),                                         //              oct.rdn
		.oct_rup                   (m2_ddr2_oct_rup),                                         //                 .rup
		.pll_mem_clk               (m2_ddr2_memory_pll_sharing_pll_mem_clk),                  //      pll_sharing.pll_mem_clk
		.pll_write_clk             (m2_ddr2_memory_pll_sharing_pll_write_clk),                //                 .pll_write_clk
		.pll_locked                (m2_ddr2_memory_pll_sharing_pll_locked),                   //                 .pll_locked
		.pll_write_clk_pre_phy_clk (m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk),    //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk),             //                 .pll_addr_cmd_clk
		.pll_avl_clk               (m2_ddr2_memory_pll_sharing_pll_avl_clk),                  //                 .pll_avl_clk
		.pll_config_clk            (m2_ddr2_memory_pll_sharing_pll_config_clk),               //                 .pll_config_clk
		.dll_pll_locked            (m2_ddr2_memory_dll_sharing_dll_pll_locked),               //      dll_sharing.dll_pll_locked
		.dll_delayctrl             (m2_ddr2_memory_dll_sharing_dll_delayctrl)                 //                 .dll_delayctrl
	);

	MebX_Qsys_Project_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (m2_ddr2_memory_afi_half_clk_clk),                            //                       clk.clk
		.reset_n                             (~rst_controller_022_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_022_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_burstcount                        (nios2_gen2_0_instruction_master_burstcount),                 //                          .burstcount
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	MebX_Qsys_Project_onchip_memory onchip_memory (
		.clk        (m2_ddr2_memory_afi_half_clk_clk),               //   clk1.clk
		.address    (mm_interconnect_1_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_1_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_008_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_008_reset_out_reset_req),        //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	MebX_Qsys_Project_pio_BUTTON pio_button (
		.clk      (clk50_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_019_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_2_pio_button_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_pio_button_s1_readdata), //                    .readdata
		.in_port  (button_export)                             // external_connection.export
	);

	MebX_Qsys_Project_pio_DIP pio_dip (
		.clk      (clk50_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_019_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_2_pio_dip_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_pio_dip_s1_readdata), //                    .readdata
		.in_port  (dip_export)                             // external_connection.export
	);

	MebX_Qsys_Project_pio_EXT pio_ext (
		.clk      (clk50_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_019_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_2_pio_ext_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_pio_ext_s1_readdata), //                    .readdata
		.in_port  (ext_export)                             // external_connection.export
	);

	MebX_Qsys_Project_pio_LED pio_led (
		.clk        (clk50_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_2_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_pio_led_s1_readdata),   //                    .readdata
		.out_port   (led_de4_export)                           // external_connection.export
	);

	MebX_Qsys_Project_pio_LED_painel pio_led_painel (
		.clk        (clk50_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_2_pio_led_painel_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_pio_led_painel_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_pio_led_painel_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_pio_led_painel_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_pio_led_painel_s1_readdata),   //                    .readdata
		.out_port   (led_painel_export)                               // external_connection.export
	);

	MebX_Qsys_Project_pio_ctrl_io_lvds pio_ctrl_io_lvds (
		.clk        (clk50_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_2_pio_ctrl_io_lvds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_pio_ctrl_io_lvds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_pio_ctrl_io_lvds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_pio_ctrl_io_lvds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_pio_ctrl_io_lvds_s1_readdata),   //                    .readdata
		.out_port   (ctrl_io_lvds_export)                               // external_connection.export
	);

	nrme_rmap_memory_nfee_area_top rmap_mem_nfee_comm_1 (
		.reset_i                             (rst_controller_002_reset_out_reset),                                                //                      reset_sink.reset
		.clk_100_i                           (m2_ddr2_memory_afi_half_clk_clk),                                                   //               clock_sink_100mhz.clk
		.avs_0_rmap_address_i                (mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_address),                //             avalon_rmap_slave_0.address
		.avs_0_rmap_write_i                  (mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_write),                  //                                .write
		.avs_0_rmap_read_i                   (mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_read),                   //                                .read
		.avs_0_rmap_readdata_o               (mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_readdata),               //                                .readdata
		.avs_0_rmap_writedata_i              (mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_writedata),              //                                .writedata
		.avs_0_rmap_waitrequest_o            (mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_waitrequest),            //                                .waitrequest
		.avs_0_rmap_byteenable_i             (mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_byteenable),             //                                .byteenable
		.fee_0_rmap_wr_address_i             (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_wr_address_signal),         //    conduit_end_fee_rmap_slave_0.wr_address_signal
		.fee_0_rmap_write_i                  (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_write_signal),              //                                .write_signal
		.fee_0_rmap_writedata_i              (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_writedata_signal),          //                                .writedata_signal
		.fee_0_rmap_rd_address_i             (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_rd_address_signal),         //                                .rd_address_signal
		.fee_0_rmap_read_i                   (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_codec_read_signal),               //                                .read_signal
		.fee_0_rmap_wr_waitrequest_o         (rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal),           //                                .wr_waitrequest_signal
		.fee_0_rmap_readdata_o               (rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_readdata_signal),                 //                                .readdata_signal
		.fee_0_rmap_rd_waitrequest_o         (rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal),           //                                .rd_waitrequest_signal
		.fee_1_rmap_wr_address_i             (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_wr_address_signal),            //    conduit_end_fee_rmap_slave_1.wr_address_signal
		.fee_1_rmap_write_i                  (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_write_signal),                 //                                .write_signal
		.fee_1_rmap_writedata_i              (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_writedata_signal),             //                                .writedata_signal
		.fee_1_rmap_rd_address_i             (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_rd_address_signal),            //                                .rd_address_signal
		.fee_1_rmap_read_i                   (comm_pedreiro_v1_01_1_conduit_end_fee_rmap_master_hk_read_signal),                  //                                .read_signal
		.fee_1_rmap_wr_waitrequest_o         (rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal),           //                                .wr_waitrequest_signal
		.fee_1_rmap_readdata_o               (rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_readdata_signal),                 //                                .readdata_signal
		.fee_1_rmap_rd_waitrequest_o         (rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal),           //                                .rd_waitrequest_signal
		.channel_hk_timecode_control_i       (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_timecode_control_signal),          //       conduit_end_channel_hk_in.timecode_control_signal
		.channel_hk_timecode_time_i          (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_timecode_time_signal),             //                                .timecode_time_signal
		.channel_hk_rmap_target_status_i     (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_rmap_target_status_signal),        //                                .rmap_target_status_signal
		.channel_hk_rmap_target_indicate_i   (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_rmap_target_indicate_signal),      //                                .rmap_target_indicate_signal
		.channel_hk_spw_link_escape_err_i    (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_escape_err_signal),       //                                .spw_link_escape_err_signal
		.channel_hk_spw_link_credit_err_i    (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_credit_err_signal),       //                                .spw_link_credit_err_signal
		.channel_hk_spw_link_parity_err_i    (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_parity_err_signal),       //                                .spw_link_parity_err_signal
		.channel_hk_spw_link_disconnect_i    (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_disconnect_signal),       //                                .spw_link_disconnect_signal
		.channel_hk_spw_link_running_i       (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_spw_link_running_signal),          //                                .spw_link_running_signal
		.channel_hk_frame_counter_i          (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_frame_counter_signal),             //                                .frame_counter_signal
		.channel_hk_frame_number_i           (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_frame_number_signal),              //                                .frame_number_signal
		.channel_hk_err_win_wrong_x_coord_i  (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal),     //                                .err_win_wrong_x_coord_signal
		.channel_hk_err_win_wrong_y_coord_i  (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal),     //                                .err_win_wrong_y_coord_signal
		.channel_hk_err_e_side_buffer_full_i (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_e_side_buffer_full_signal),    //                                .err_e_side_buffer_full_signal
		.channel_hk_err_f_side_buffer_full_i (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_f_side_buffer_full_signal),    //                                .err_f_side_buffer_full_signal
		.channel_hk_err_invalid_ccd_mode_i   (comm_pedreiro_v1_01_1_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal),      //                                .err_invalid_ccd_mode_signal
		.avm_rmap_readdata_i                 (rmap_mem_nfee_comm_1_avalon_mm_rmap_master_readdata),                               //           avalon_mm_rmap_master.readdata
		.avm_rmap_waitrequest_i              (rmap_mem_nfee_comm_1_avalon_mm_rmap_master_waitrequest),                            //                                .waitrequest
		.avm_rmap_address_o                  (rmap_mem_nfee_comm_1_avalon_mm_rmap_master_address),                                //                                .address
		.avm_rmap_read_o                     (rmap_mem_nfee_comm_1_avalon_mm_rmap_master_read),                                   //                                .read
		.avm_rmap_write_o                    (rmap_mem_nfee_comm_1_avalon_mm_rmap_master_write),                                  //                                .write
		.avm_rmap_writedata_o                (rmap_mem_nfee_comm_1_avalon_mm_rmap_master_writedata),                              //                                .writedata
		.channel_win_mem_addr_offset_i       (comm_pedreiro_v1_01_1_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal)  // conduit_end_rmap_avm_configs_in.win_mem_addr_offset_signal
	);

	nrme_rmap_memory_nfee_area_top rmap_mem_nfee_comm_2 (
		.reset_i                             (rst_controller_003_reset_out_reset),                                                //                      reset_sink.reset
		.clk_100_i                           (m2_ddr2_memory_afi_half_clk_clk),                                                   //               clock_sink_100mhz.clk
		.avs_0_rmap_address_i                (mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_address),                //             avalon_rmap_slave_0.address
		.avs_0_rmap_write_i                  (mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_write),                  //                                .write
		.avs_0_rmap_read_i                   (mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_read),                   //                                .read
		.avs_0_rmap_readdata_o               (mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_readdata),               //                                .readdata
		.avs_0_rmap_writedata_i              (mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_writedata),              //                                .writedata
		.avs_0_rmap_waitrequest_o            (mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_waitrequest),            //                                .waitrequest
		.avs_0_rmap_byteenable_i             (mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_byteenable),             //                                .byteenable
		.fee_0_rmap_wr_address_i             (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_wr_address_signal),         //    conduit_end_fee_rmap_slave_0.wr_address_signal
		.fee_0_rmap_write_i                  (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_write_signal),              //                                .write_signal
		.fee_0_rmap_writedata_i              (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_writedata_signal),          //                                .writedata_signal
		.fee_0_rmap_rd_address_i             (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_rd_address_signal),         //                                .rd_address_signal
		.fee_0_rmap_read_i                   (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_codec_read_signal),               //                                .read_signal
		.fee_0_rmap_wr_waitrequest_o         (rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal),           //                                .wr_waitrequest_signal
		.fee_0_rmap_readdata_o               (rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_readdata_signal),                 //                                .readdata_signal
		.fee_0_rmap_rd_waitrequest_o         (rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal),           //                                .rd_waitrequest_signal
		.fee_1_rmap_wr_address_i             (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_wr_address_signal),            //    conduit_end_fee_rmap_slave_1.wr_address_signal
		.fee_1_rmap_write_i                  (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_write_signal),                 //                                .write_signal
		.fee_1_rmap_writedata_i              (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_writedata_signal),             //                                .writedata_signal
		.fee_1_rmap_rd_address_i             (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_rd_address_signal),            //                                .rd_address_signal
		.fee_1_rmap_read_i                   (comm_pedreiro_v1_01_2_conduit_end_fee_rmap_master_hk_read_signal),                  //                                .read_signal
		.fee_1_rmap_wr_waitrequest_o         (rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal),           //                                .wr_waitrequest_signal
		.fee_1_rmap_readdata_o               (rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_readdata_signal),                 //                                .readdata_signal
		.fee_1_rmap_rd_waitrequest_o         (rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal),           //                                .rd_waitrequest_signal
		.channel_hk_timecode_control_i       (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_timecode_control_signal),          //       conduit_end_channel_hk_in.timecode_control_signal
		.channel_hk_timecode_time_i          (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_timecode_time_signal),             //                                .timecode_time_signal
		.channel_hk_rmap_target_status_i     (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_rmap_target_status_signal),        //                                .rmap_target_status_signal
		.channel_hk_rmap_target_indicate_i   (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_rmap_target_indicate_signal),      //                                .rmap_target_indicate_signal
		.channel_hk_spw_link_escape_err_i    (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_escape_err_signal),       //                                .spw_link_escape_err_signal
		.channel_hk_spw_link_credit_err_i    (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_credit_err_signal),       //                                .spw_link_credit_err_signal
		.channel_hk_spw_link_parity_err_i    (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_parity_err_signal),       //                                .spw_link_parity_err_signal
		.channel_hk_spw_link_disconnect_i    (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_disconnect_signal),       //                                .spw_link_disconnect_signal
		.channel_hk_spw_link_running_i       (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_spw_link_running_signal),          //                                .spw_link_running_signal
		.channel_hk_frame_counter_i          (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_frame_counter_signal),             //                                .frame_counter_signal
		.channel_hk_frame_number_i           (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_frame_number_signal),              //                                .frame_number_signal
		.channel_hk_err_win_wrong_x_coord_i  (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal),     //                                .err_win_wrong_x_coord_signal
		.channel_hk_err_win_wrong_y_coord_i  (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal),     //                                .err_win_wrong_y_coord_signal
		.channel_hk_err_e_side_buffer_full_i (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_e_side_buffer_full_signal),    //                                .err_e_side_buffer_full_signal
		.channel_hk_err_f_side_buffer_full_i (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_f_side_buffer_full_signal),    //                                .err_f_side_buffer_full_signal
		.channel_hk_err_invalid_ccd_mode_i   (comm_pedreiro_v1_01_2_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal),      //                                .err_invalid_ccd_mode_signal
		.avm_rmap_readdata_i                 (rmap_mem_nfee_comm_2_avalon_mm_rmap_master_readdata),                               //           avalon_mm_rmap_master.readdata
		.avm_rmap_waitrequest_i              (rmap_mem_nfee_comm_2_avalon_mm_rmap_master_waitrequest),                            //                                .waitrequest
		.avm_rmap_address_o                  (rmap_mem_nfee_comm_2_avalon_mm_rmap_master_address),                                //                                .address
		.avm_rmap_read_o                     (rmap_mem_nfee_comm_2_avalon_mm_rmap_master_read),                                   //                                .read
		.avm_rmap_write_o                    (rmap_mem_nfee_comm_2_avalon_mm_rmap_master_write),                                  //                                .write
		.avm_rmap_writedata_o                (rmap_mem_nfee_comm_2_avalon_mm_rmap_master_writedata),                              //                                .writedata
		.channel_win_mem_addr_offset_i       (comm_pedreiro_v1_01_2_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal)  // conduit_end_rmap_avm_configs_in.win_mem_addr_offset_signal
	);

	nrme_rmap_memory_nfee_area_top rmap_mem_nfee_comm_3 (
		.reset_i                             (rst_controller_004_reset_out_reset),                                                //                      reset_sink.reset
		.clk_100_i                           (m2_ddr2_memory_afi_half_clk_clk),                                                   //               clock_sink_100mhz.clk
		.avs_0_rmap_address_i                (mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_address),                //             avalon_rmap_slave_0.address
		.avs_0_rmap_write_i                  (mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_write),                  //                                .write
		.avs_0_rmap_read_i                   (mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_read),                   //                                .read
		.avs_0_rmap_readdata_o               (mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_readdata),               //                                .readdata
		.avs_0_rmap_writedata_i              (mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_writedata),              //                                .writedata
		.avs_0_rmap_waitrequest_o            (mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_waitrequest),            //                                .waitrequest
		.avs_0_rmap_byteenable_i             (mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_byteenable),             //                                .byteenable
		.fee_0_rmap_wr_address_i             (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_wr_address_signal),         //    conduit_end_fee_rmap_slave_0.wr_address_signal
		.fee_0_rmap_write_i                  (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_write_signal),              //                                .write_signal
		.fee_0_rmap_writedata_i              (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_writedata_signal),          //                                .writedata_signal
		.fee_0_rmap_rd_address_i             (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_rd_address_signal),         //                                .rd_address_signal
		.fee_0_rmap_read_i                   (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_codec_read_signal),               //                                .read_signal
		.fee_0_rmap_wr_waitrequest_o         (rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal),           //                                .wr_waitrequest_signal
		.fee_0_rmap_readdata_o               (rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_readdata_signal),                 //                                .readdata_signal
		.fee_0_rmap_rd_waitrequest_o         (rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal),           //                                .rd_waitrequest_signal
		.fee_1_rmap_wr_address_i             (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_wr_address_signal),            //    conduit_end_fee_rmap_slave_1.wr_address_signal
		.fee_1_rmap_write_i                  (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_write_signal),                 //                                .write_signal
		.fee_1_rmap_writedata_i              (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_writedata_signal),             //                                .writedata_signal
		.fee_1_rmap_rd_address_i             (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_rd_address_signal),            //                                .rd_address_signal
		.fee_1_rmap_read_i                   (comm_pedreiro_v1_01_3_conduit_end_fee_rmap_master_hk_read_signal),                  //                                .read_signal
		.fee_1_rmap_wr_waitrequest_o         (rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal),           //                                .wr_waitrequest_signal
		.fee_1_rmap_readdata_o               (rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_readdata_signal),                 //                                .readdata_signal
		.fee_1_rmap_rd_waitrequest_o         (rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal),           //                                .rd_waitrequest_signal
		.channel_hk_timecode_control_i       (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_timecode_control_signal),          //       conduit_end_channel_hk_in.timecode_control_signal
		.channel_hk_timecode_time_i          (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_timecode_time_signal),             //                                .timecode_time_signal
		.channel_hk_rmap_target_status_i     (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_rmap_target_status_signal),        //                                .rmap_target_status_signal
		.channel_hk_rmap_target_indicate_i   (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_rmap_target_indicate_signal),      //                                .rmap_target_indicate_signal
		.channel_hk_spw_link_escape_err_i    (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_escape_err_signal),       //                                .spw_link_escape_err_signal
		.channel_hk_spw_link_credit_err_i    (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_credit_err_signal),       //                                .spw_link_credit_err_signal
		.channel_hk_spw_link_parity_err_i    (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_parity_err_signal),       //                                .spw_link_parity_err_signal
		.channel_hk_spw_link_disconnect_i    (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_disconnect_signal),       //                                .spw_link_disconnect_signal
		.channel_hk_spw_link_running_i       (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_spw_link_running_signal),          //                                .spw_link_running_signal
		.channel_hk_frame_counter_i          (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_frame_counter_signal),             //                                .frame_counter_signal
		.channel_hk_frame_number_i           (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_frame_number_signal),              //                                .frame_number_signal
		.channel_hk_err_win_wrong_x_coord_i  (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal),     //                                .err_win_wrong_x_coord_signal
		.channel_hk_err_win_wrong_y_coord_i  (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal),     //                                .err_win_wrong_y_coord_signal
		.channel_hk_err_e_side_buffer_full_i (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_e_side_buffer_full_signal),    //                                .err_e_side_buffer_full_signal
		.channel_hk_err_f_side_buffer_full_i (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_f_side_buffer_full_signal),    //                                .err_f_side_buffer_full_signal
		.channel_hk_err_invalid_ccd_mode_i   (comm_pedreiro_v1_01_3_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal),      //                                .err_invalid_ccd_mode_signal
		.avm_rmap_readdata_i                 (rmap_mem_nfee_comm_3_avalon_mm_rmap_master_readdata),                               //           avalon_mm_rmap_master.readdata
		.avm_rmap_waitrequest_i              (rmap_mem_nfee_comm_3_avalon_mm_rmap_master_waitrequest),                            //                                .waitrequest
		.avm_rmap_address_o                  (rmap_mem_nfee_comm_3_avalon_mm_rmap_master_address),                                //                                .address
		.avm_rmap_read_o                     (rmap_mem_nfee_comm_3_avalon_mm_rmap_master_read),                                   //                                .read
		.avm_rmap_write_o                    (rmap_mem_nfee_comm_3_avalon_mm_rmap_master_write),                                  //                                .write
		.avm_rmap_writedata_o                (rmap_mem_nfee_comm_3_avalon_mm_rmap_master_writedata),                              //                                .writedata
		.channel_win_mem_addr_offset_i       (comm_pedreiro_v1_01_3_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal)  // conduit_end_rmap_avm_configs_in.win_mem_addr_offset_signal
	);

	nrme_rmap_memory_nfee_area_top rmap_mem_nfee_comm_4 (
		.reset_i                             (rst_controller_005_reset_out_reset),                                                //                      reset_sink.reset
		.clk_100_i                           (m2_ddr2_memory_afi_half_clk_clk),                                                   //               clock_sink_100mhz.clk
		.avs_0_rmap_address_i                (mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_address),                //             avalon_rmap_slave_0.address
		.avs_0_rmap_write_i                  (mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_write),                  //                                .write
		.avs_0_rmap_read_i                   (mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_read),                   //                                .read
		.avs_0_rmap_readdata_o               (mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_readdata),               //                                .readdata
		.avs_0_rmap_writedata_i              (mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_writedata),              //                                .writedata
		.avs_0_rmap_waitrequest_o            (mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_waitrequest),            //                                .waitrequest
		.avs_0_rmap_byteenable_i             (mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_byteenable),             //                                .byteenable
		.fee_0_rmap_wr_address_i             (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_wr_address_signal),         //    conduit_end_fee_rmap_slave_0.wr_address_signal
		.fee_0_rmap_write_i                  (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_write_signal),              //                                .write_signal
		.fee_0_rmap_writedata_i              (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_writedata_signal),          //                                .writedata_signal
		.fee_0_rmap_rd_address_i             (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_rd_address_signal),         //                                .rd_address_signal
		.fee_0_rmap_read_i                   (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_codec_read_signal),               //                                .read_signal
		.fee_0_rmap_wr_waitrequest_o         (rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal),           //                                .wr_waitrequest_signal
		.fee_0_rmap_readdata_o               (rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_readdata_signal),                 //                                .readdata_signal
		.fee_0_rmap_rd_waitrequest_o         (rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal),           //                                .rd_waitrequest_signal
		.fee_1_rmap_wr_address_i             (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_wr_address_signal),            //    conduit_end_fee_rmap_slave_1.wr_address_signal
		.fee_1_rmap_write_i                  (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_write_signal),                 //                                .write_signal
		.fee_1_rmap_writedata_i              (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_writedata_signal),             //                                .writedata_signal
		.fee_1_rmap_rd_address_i             (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_rd_address_signal),            //                                .rd_address_signal
		.fee_1_rmap_read_i                   (comm_pedreiro_v1_01_4_conduit_end_fee_rmap_master_hk_read_signal),                  //                                .read_signal
		.fee_1_rmap_wr_waitrequest_o         (rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal),           //                                .wr_waitrequest_signal
		.fee_1_rmap_readdata_o               (rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_readdata_signal),                 //                                .readdata_signal
		.fee_1_rmap_rd_waitrequest_o         (rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal),           //                                .rd_waitrequest_signal
		.channel_hk_timecode_control_i       (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_timecode_control_signal),          //       conduit_end_channel_hk_in.timecode_control_signal
		.channel_hk_timecode_time_i          (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_timecode_time_signal),             //                                .timecode_time_signal
		.channel_hk_rmap_target_status_i     (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_rmap_target_status_signal),        //                                .rmap_target_status_signal
		.channel_hk_rmap_target_indicate_i   (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_rmap_target_indicate_signal),      //                                .rmap_target_indicate_signal
		.channel_hk_spw_link_escape_err_i    (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_escape_err_signal),       //                                .spw_link_escape_err_signal
		.channel_hk_spw_link_credit_err_i    (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_credit_err_signal),       //                                .spw_link_credit_err_signal
		.channel_hk_spw_link_parity_err_i    (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_parity_err_signal),       //                                .spw_link_parity_err_signal
		.channel_hk_spw_link_disconnect_i    (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_disconnect_signal),       //                                .spw_link_disconnect_signal
		.channel_hk_spw_link_running_i       (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_spw_link_running_signal),          //                                .spw_link_running_signal
		.channel_hk_frame_counter_i          (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_frame_counter_signal),             //                                .frame_counter_signal
		.channel_hk_frame_number_i           (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_frame_number_signal),              //                                .frame_number_signal
		.channel_hk_err_win_wrong_x_coord_i  (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal),     //                                .err_win_wrong_x_coord_signal
		.channel_hk_err_win_wrong_y_coord_i  (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal),     //                                .err_win_wrong_y_coord_signal
		.channel_hk_err_e_side_buffer_full_i (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_e_side_buffer_full_signal),    //                                .err_e_side_buffer_full_signal
		.channel_hk_err_f_side_buffer_full_i (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_f_side_buffer_full_signal),    //                                .err_f_side_buffer_full_signal
		.channel_hk_err_invalid_ccd_mode_i   (comm_pedreiro_v1_01_4_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal),      //                                .err_invalid_ccd_mode_signal
		.avm_rmap_readdata_i                 (rmap_mem_nfee_comm_4_avalon_mm_rmap_master_readdata),                               //           avalon_mm_rmap_master.readdata
		.avm_rmap_waitrequest_i              (rmap_mem_nfee_comm_4_avalon_mm_rmap_master_waitrequest),                            //                                .waitrequest
		.avm_rmap_address_o                  (rmap_mem_nfee_comm_4_avalon_mm_rmap_master_address),                                //                                .address
		.avm_rmap_read_o                     (rmap_mem_nfee_comm_4_avalon_mm_rmap_master_read),                                   //                                .read
		.avm_rmap_write_o                    (rmap_mem_nfee_comm_4_avalon_mm_rmap_master_write),                                  //                                .write
		.avm_rmap_writedata_o                (rmap_mem_nfee_comm_4_avalon_mm_rmap_master_writedata),                              //                                .writedata
		.channel_win_mem_addr_offset_i       (comm_pedreiro_v1_01_4_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal)  // conduit_end_rmap_avm_configs_in.win_mem_addr_offset_signal
	);

	nrme_rmap_memory_nfee_area_top rmap_mem_nfee_comm_5 (
		.reset_i                             (rst_controller_006_reset_out_reset),                                                //                      reset_sink.reset
		.clk_100_i                           (m2_ddr2_memory_afi_half_clk_clk),                                                   //               clock_sink_100mhz.clk
		.avs_0_rmap_address_i                (mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_address),                //             avalon_rmap_slave_0.address
		.avs_0_rmap_write_i                  (mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_write),                  //                                .write
		.avs_0_rmap_read_i                   (mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_read),                   //                                .read
		.avs_0_rmap_readdata_o               (mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_readdata),               //                                .readdata
		.avs_0_rmap_writedata_i              (mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_writedata),              //                                .writedata
		.avs_0_rmap_waitrequest_o            (mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_waitrequest),            //                                .waitrequest
		.avs_0_rmap_byteenable_i             (mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_byteenable),             //                                .byteenable
		.fee_0_rmap_wr_address_i             (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_wr_address_signal),         //    conduit_end_fee_rmap_slave_0.wr_address_signal
		.fee_0_rmap_write_i                  (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_write_signal),              //                                .write_signal
		.fee_0_rmap_writedata_i              (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_writedata_signal),          //                                .writedata_signal
		.fee_0_rmap_rd_address_i             (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_rd_address_signal),         //                                .rd_address_signal
		.fee_0_rmap_read_i                   (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_codec_read_signal),               //                                .read_signal
		.fee_0_rmap_wr_waitrequest_o         (rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal),           //                                .wr_waitrequest_signal
		.fee_0_rmap_readdata_o               (rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_readdata_signal),                 //                                .readdata_signal
		.fee_0_rmap_rd_waitrequest_o         (rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal),           //                                .rd_waitrequest_signal
		.fee_1_rmap_wr_address_i             (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_wr_address_signal),            //    conduit_end_fee_rmap_slave_1.wr_address_signal
		.fee_1_rmap_write_i                  (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_write_signal),                 //                                .write_signal
		.fee_1_rmap_writedata_i              (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_writedata_signal),             //                                .writedata_signal
		.fee_1_rmap_rd_address_i             (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_rd_address_signal),            //                                .rd_address_signal
		.fee_1_rmap_read_i                   (comm_pedreiro_v1_01_5_conduit_end_fee_rmap_master_hk_read_signal),                  //                                .read_signal
		.fee_1_rmap_wr_waitrequest_o         (rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal),           //                                .wr_waitrequest_signal
		.fee_1_rmap_readdata_o               (rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_readdata_signal),                 //                                .readdata_signal
		.fee_1_rmap_rd_waitrequest_o         (rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal),           //                                .rd_waitrequest_signal
		.channel_hk_timecode_control_i       (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_timecode_control_signal),          //       conduit_end_channel_hk_in.timecode_control_signal
		.channel_hk_timecode_time_i          (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_timecode_time_signal),             //                                .timecode_time_signal
		.channel_hk_rmap_target_status_i     (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_rmap_target_status_signal),        //                                .rmap_target_status_signal
		.channel_hk_rmap_target_indicate_i   (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_rmap_target_indicate_signal),      //                                .rmap_target_indicate_signal
		.channel_hk_spw_link_escape_err_i    (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_escape_err_signal),       //                                .spw_link_escape_err_signal
		.channel_hk_spw_link_credit_err_i    (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_credit_err_signal),       //                                .spw_link_credit_err_signal
		.channel_hk_spw_link_parity_err_i    (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_parity_err_signal),       //                                .spw_link_parity_err_signal
		.channel_hk_spw_link_disconnect_i    (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_disconnect_signal),       //                                .spw_link_disconnect_signal
		.channel_hk_spw_link_running_i       (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_spw_link_running_signal),          //                                .spw_link_running_signal
		.channel_hk_frame_counter_i          (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_frame_counter_signal),             //                                .frame_counter_signal
		.channel_hk_frame_number_i           (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_frame_number_signal),              //                                .frame_number_signal
		.channel_hk_err_win_wrong_x_coord_i  (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal),     //                                .err_win_wrong_x_coord_signal
		.channel_hk_err_win_wrong_y_coord_i  (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal),     //                                .err_win_wrong_y_coord_signal
		.channel_hk_err_e_side_buffer_full_i (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_e_side_buffer_full_signal),    //                                .err_e_side_buffer_full_signal
		.channel_hk_err_f_side_buffer_full_i (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_f_side_buffer_full_signal),    //                                .err_f_side_buffer_full_signal
		.channel_hk_err_invalid_ccd_mode_i   (comm_pedreiro_v1_01_5_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal),      //                                .err_invalid_ccd_mode_signal
		.avm_rmap_readdata_i                 (rmap_mem_nfee_comm_5_avalon_mm_rmap_master_readdata),                               //           avalon_mm_rmap_master.readdata
		.avm_rmap_waitrequest_i              (rmap_mem_nfee_comm_5_avalon_mm_rmap_master_waitrequest),                            //                                .waitrequest
		.avm_rmap_address_o                  (rmap_mem_nfee_comm_5_avalon_mm_rmap_master_address),                                //                                .address
		.avm_rmap_read_o                     (rmap_mem_nfee_comm_5_avalon_mm_rmap_master_read),                                   //                                .read
		.avm_rmap_write_o                    (rmap_mem_nfee_comm_5_avalon_mm_rmap_master_write),                                  //                                .write
		.avm_rmap_writedata_o                (rmap_mem_nfee_comm_5_avalon_mm_rmap_master_writedata),                              //                                .writedata
		.channel_win_mem_addr_offset_i       (comm_pedreiro_v1_01_5_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal)  // conduit_end_rmap_avm_configs_in.win_mem_addr_offset_signal
	);

	nrme_rmap_memory_nfee_area_top rmap_mem_nfee_comm_6 (
		.reset_i                             (rst_controller_007_reset_out_reset),                                                //                      reset_sink.reset
		.clk_100_i                           (m2_ddr2_memory_afi_half_clk_clk),                                                   //               clock_sink_100mhz.clk
		.avs_0_rmap_address_i                (mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_address),                //             avalon_rmap_slave_0.address
		.avs_0_rmap_write_i                  (mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_write),                  //                                .write
		.avs_0_rmap_read_i                   (mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_read),                   //                                .read
		.avs_0_rmap_readdata_o               (mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_readdata),               //                                .readdata
		.avs_0_rmap_writedata_i              (mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_writedata),              //                                .writedata
		.avs_0_rmap_waitrequest_o            (mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_waitrequest),            //                                .waitrequest
		.avs_0_rmap_byteenable_i             (mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_byteenable),             //                                .byteenable
		.fee_0_rmap_wr_address_i             (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_wr_address_signal),         //    conduit_end_fee_rmap_slave_0.wr_address_signal
		.fee_0_rmap_write_i                  (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_write_signal),              //                                .write_signal
		.fee_0_rmap_writedata_i              (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_writedata_signal),          //                                .writedata_signal
		.fee_0_rmap_rd_address_i             (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_rd_address_signal),         //                                .rd_address_signal
		.fee_0_rmap_read_i                   (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_codec_read_signal),               //                                .read_signal
		.fee_0_rmap_wr_waitrequest_o         (rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal),           //                                .wr_waitrequest_signal
		.fee_0_rmap_readdata_o               (rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_readdata_signal),                 //                                .readdata_signal
		.fee_0_rmap_rd_waitrequest_o         (rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal),           //                                .rd_waitrequest_signal
		.fee_1_rmap_wr_address_i             (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_wr_address_signal),            //    conduit_end_fee_rmap_slave_1.wr_address_signal
		.fee_1_rmap_write_i                  (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_write_signal),                 //                                .write_signal
		.fee_1_rmap_writedata_i              (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_writedata_signal),             //                                .writedata_signal
		.fee_1_rmap_rd_address_i             (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_rd_address_signal),            //                                .rd_address_signal
		.fee_1_rmap_read_i                   (comm_pedreiro_v1_01_6_conduit_end_fee_rmap_master_hk_read_signal),                  //                                .read_signal
		.fee_1_rmap_wr_waitrequest_o         (rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal),           //                                .wr_waitrequest_signal
		.fee_1_rmap_readdata_o               (rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_readdata_signal),                 //                                .readdata_signal
		.fee_1_rmap_rd_waitrequest_o         (rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal),           //                                .rd_waitrequest_signal
		.channel_hk_timecode_control_i       (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_timecode_control_signal),          //       conduit_end_channel_hk_in.timecode_control_signal
		.channel_hk_timecode_time_i          (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_timecode_time_signal),             //                                .timecode_time_signal
		.channel_hk_rmap_target_status_i     (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_rmap_target_status_signal),        //                                .rmap_target_status_signal
		.channel_hk_rmap_target_indicate_i   (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_rmap_target_indicate_signal),      //                                .rmap_target_indicate_signal
		.channel_hk_spw_link_escape_err_i    (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_escape_err_signal),       //                                .spw_link_escape_err_signal
		.channel_hk_spw_link_credit_err_i    (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_credit_err_signal),       //                                .spw_link_credit_err_signal
		.channel_hk_spw_link_parity_err_i    (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_parity_err_signal),       //                                .spw_link_parity_err_signal
		.channel_hk_spw_link_disconnect_i    (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_disconnect_signal),       //                                .spw_link_disconnect_signal
		.channel_hk_spw_link_running_i       (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_spw_link_running_signal),          //                                .spw_link_running_signal
		.channel_hk_frame_counter_i          (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_frame_counter_signal),             //                                .frame_counter_signal
		.channel_hk_frame_number_i           (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_frame_number_signal),              //                                .frame_number_signal
		.channel_hk_err_win_wrong_x_coord_i  (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_win_wrong_x_coord_signal),     //                                .err_win_wrong_x_coord_signal
		.channel_hk_err_win_wrong_y_coord_i  (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_win_wrong_y_coord_signal),     //                                .err_win_wrong_y_coord_signal
		.channel_hk_err_e_side_buffer_full_i (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_e_side_buffer_full_signal),    //                                .err_e_side_buffer_full_signal
		.channel_hk_err_f_side_buffer_full_i (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_f_side_buffer_full_signal),    //                                .err_f_side_buffer_full_signal
		.channel_hk_err_invalid_ccd_mode_i   (comm_pedreiro_v1_01_6_conduit_end_channel_hk_out_err_invalid_ccd_mode_signal),      //                                .err_invalid_ccd_mode_signal
		.avm_rmap_readdata_i                 (rmap_mem_nfee_comm_6_avalon_mm_rmap_master_readdata),                               //           avalon_mm_rmap_master.readdata
		.avm_rmap_waitrequest_i              (rmap_mem_nfee_comm_6_avalon_mm_rmap_master_waitrequest),                            //                                .waitrequest
		.avm_rmap_address_o                  (rmap_mem_nfee_comm_6_avalon_mm_rmap_master_address),                                //                                .address
		.avm_rmap_read_o                     (rmap_mem_nfee_comm_6_avalon_mm_rmap_master_read),                                   //                                .read
		.avm_rmap_write_o                    (rmap_mem_nfee_comm_6_avalon_mm_rmap_master_write),                                  //                                .write
		.avm_rmap_writedata_o                (rmap_mem_nfee_comm_6_avalon_mm_rmap_master_writedata),                              //                                .writedata
		.channel_win_mem_addr_offset_i       (comm_pedreiro_v1_01_6_conduit_end_rmap_avm_configs_out_win_mem_addr_offset_signal)  // conduit_end_rmap_avm_configs_in.win_mem_addr_offset_signal
	);

	MebX_Qsys_Project_rs232_uart rs232_uart (
		.clk           (clk50_clk),                                     //                 clk.clk
		.reset_n       (~rst_controller_023_reset_out_reset),           //               reset.reset_n
		.address       (mm_interconnect_2_rs232_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_2_rs232_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_2_rs232_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_2_rs232_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_2_rs232_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_2_rs232_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_2_rs232_uart_s1_readdata),      //                    .readdata
		.rxd           (rs232_uart_rxd),                                // external_connection.export
		.txd           (rs232_uart_txd),                                //                    .export
		.irq           (irq_synchronizer_002_receiver_irq)              //                 irq.irq
	);

	rst_controller_top rst_controller (
		.clock_sink_clk                          (clk50_clk),                                                                //                  clock_sink.clk
		.reset_sink_reset                        (rst_controller_019_reset_out_reset),                                       //                  reset_sink.reset
		.reset_source_ftdi_reset                 (),                                                                         //           reset_source_ftdi.reset
		.reset_source_sync_reset                 (rst_controller_reset_source_sync_reset),                                   //           reset_source_sync.reset
		.reset_source_rs232_reset                (rst_controller_reset_source_rs232_reset),                                  //          reset_source_rs232.reset
		.reset_source_sd_card_reset              (rst_controller_reset_source_sd_card_reset),                                //        reset_source_sd_card.reset
		.reset_source_comm_ch8_reset             (rst_controller_reset_source_comm_ch8_reset),                               //       reset_source_comm_ch8.reset
		.reset_source_comm_ch7_reset             (rst_controller_reset_source_comm_ch7_reset),                               //       reset_source_comm_ch7.reset
		.reset_source_comm_ch6_reset             (rst_controller_reset_source_comm_ch6_reset),                               //       reset_source_comm_ch6.reset
		.reset_source_comm_ch5_reset             (rst_controller_reset_source_comm_ch5_reset),                               //       reset_source_comm_ch5.reset
		.reset_source_comm_ch4_reset             (rst_controller_reset_source_comm_ch4_reset),                               //       reset_source_comm_ch4.reset
		.reset_source_comm_ch3_reset             (rst_controller_reset_source_comm_ch3_reset),                               //       reset_source_comm_ch3.reset
		.reset_source_comm_ch2_reset             (rst_controller_reset_source_comm_ch2_reset),                               //       reset_source_comm_ch2.reset
		.reset_source_comm_ch1_reset             (rst_controller_reset_source_comm_ch1_reset),                               //       reset_source_comm_ch1.reset
		.avalon_slave_rst_controller_address     (mm_interconnect_2_rst_controller_avalon_rst_controller_slave_address),     // avalon_rst_controller_slave.address
		.avalon_slave_rst_controller_write       (mm_interconnect_2_rst_controller_avalon_rst_controller_slave_write),       //                            .write
		.avalon_slave_rst_controller_read        (mm_interconnect_2_rst_controller_avalon_rst_controller_slave_read),        //                            .read
		.avalon_slave_rst_controller_writedata   (mm_interconnect_2_rst_controller_avalon_rst_controller_slave_writedata),   //                            .writedata
		.avalon_slave_rst_controller_readdata    (mm_interconnect_2_rst_controller_avalon_rst_controller_slave_readdata),    //                            .readdata
		.avalon_slave_rst_controller_waitrequest (mm_interconnect_2_rst_controller_avalon_rst_controller_slave_waitrequest), //                            .waitrequest
		.simucam_reset_signal                    (rst_controller_conduit_simucam_reset_t_simucam_reset_signal),              //       conduit_simucam_reset.t_simucam_reset_signal
		.reset_input_signal                      (rst_controller_conduit_reset_input_t_reset_input_signal)                   //         conduit_reset_input.t_reset_input_signal
	);

	MebX_Qsys_Project_csense_sdo rtcc_alarm (
		.clk      (clk50_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_019_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_2_rtcc_alarm_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_rtcc_alarm_s1_readdata), //                    .readdata
		.in_port  (rtcc_alarm_export)                         // external_connection.export
	);

	MebX_Qsys_Project_csense_adc_fo rtcc_cs_n (
		.clk        (clk50_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_2_rtcc_cs_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_rtcc_cs_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_rtcc_cs_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_rtcc_cs_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_rtcc_cs_n_s1_readdata),   //                    .readdata
		.out_port   (rtcc_cs_n_export)                           // external_connection.export
	);

	MebX_Qsys_Project_csense_adc_fo rtcc_sck (
		.clk        (clk50_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_2_rtcc_sck_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_rtcc_sck_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_rtcc_sck_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_rtcc_sck_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_rtcc_sck_s1_readdata),   //                    .readdata
		.out_port   (rtcc_sck_export)                           // external_connection.export
	);

	MebX_Qsys_Project_csense_adc_fo rtcc_sdi (
		.clk        (clk50_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_2_rtcc_sdi_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_rtcc_sdi_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_rtcc_sdi_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_rtcc_sdi_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_rtcc_sdi_s1_readdata),   //                    .readdata
		.out_port   (rtcc_sdi_export)                           // external_connection.export
	);

	MebX_Qsys_Project_csense_sdo rtcc_sdo (
		.clk      (clk50_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_019_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_2_rtcc_sdo_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_rtcc_sdo_s1_readdata), //                    .readdata
		.in_port  (rtcc_sdo_export)                         // external_connection.export
	);

	MebX_Qsys_Project_csense_sdo sd_card_wp_n (
		.clk      (clk50_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_019_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_2_sd_card_wp_n_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_sd_card_wp_n_s1_readdata), //                    .readdata
		.in_port  (sd_card_wp_n_io_export)                      // external_connection.export
	);

	sync_ent #(
		.g_SYNC_IRQ_NUMBER     (11),
		.g_PRE_SYNC_IRQ_NUMBER (12)
	) sync (
		.clock_sink_clk_i                (clk50_clk),                                          //                     clock.clk
		.reset_sink_reset_i              (rst_controller_024_reset_out_reset),                 //                     reset.reset
		.avalon_slave_address_i          (mm_interconnect_2_sync_avalon_mm_slave_address),     //           avalon_mm_slave.address
		.avalon_slave_read_i             (mm_interconnect_2_sync_avalon_mm_slave_read),        //                          .read
		.avalon_slave_write_i            (mm_interconnect_2_sync_avalon_mm_slave_write),       //                          .write
		.avalon_slave_writedata_i        (mm_interconnect_2_sync_avalon_mm_slave_writedata),   //                          .writedata
		.avalon_slave_byteenable_i       (mm_interconnect_2_sync_avalon_mm_slave_byteenable),  //                          .byteenable
		.avalon_slave_readdata_o         (mm_interconnect_2_sync_avalon_mm_slave_readdata),    //                          .readdata
		.avalon_slave_waitrequest_o      (mm_interconnect_2_sync_avalon_mm_slave_waitrequest), //                          .waitrequest
		.conduit_sync_signal_syncin_i    (sync_in_conduit),                                    //                   sync_in.conduit
		.conduit_sync_signal_spw1_o      (sync_spw1_conduit),                                  //                 sync_spw1.conduit
		.conduit_sync_signal_spw2_o      (sync_spw2_conduit),                                  //                 sync_spw2.conduit
		.conduit_sync_signal_spw3_o      (sync_spw3_conduit),                                  //                 sync_spw3.conduit
		.conduit_sync_signal_spw4_o      (sync_spw4_conduit),                                  //                 sync_spw4.conduit
		.conduit_sync_signal_spw5_o      (sync_spw5_conduit),                                  //                 sync_spw5.conduit
		.conduit_sync_signal_spw6_o      (sync_spw6_conduit),                                  //                 sync_spw6.conduit
		.conduit_sync_signal_spw7_o      (sync_spw7_conduit),                                  //                 sync_spw7.conduit
		.conduit_sync_signal_spw8_o      (sync_spw8_conduit),                                  //                 sync_spw8.conduit
		.conduit_sync_signal_syncout_o   (sync_out_conduit),                                   //                  sync_out.conduit
		.sync_interrupt_sender_irq_o     (irq_synchronizer_004_receiver_irq),                  //     sync_interrupt_sender.irq
		.pre_sync_interrupt_sender_irq_o (irq_synchronizer_003_receiver_irq)                   // pre_sync_interrupt_sender.irq
	);

	MebX_Qsys_Project_sysid_qsys sysid_qsys (
		.clock    (m2_ddr2_memory_afi_half_clk_clk),                     //           clk.clk
		.reset_n  (~rst_controller_008_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_qsys_control_slave_address)   //              .address
	);

	MebX_Qsys_Project_csense_adc_fo temp_scl (
		.clk        (clk50_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_2_temp_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_temp_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_temp_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_temp_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_temp_scl_s1_readdata),   //                    .readdata
		.out_port   (temp_scl_export)                           // external_connection.export
	);

	MebX_Qsys_Project_m1_ddr2_i2c_sda temp_sda (
		.clk        (clk50_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_019_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_2_temp_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_temp_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_temp_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_temp_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_temp_sda_s1_readdata),   //                    .readdata
		.bidir_port (temp_sda_export)                           // external_connection.export
	);

	MebX_Qsys_Project_timer_1ms timer_1ms (
		.clk           (clk50_clk),                                 //           clk.clk
		.reset_n       (~rst_controller_019_reset_out_reset),       //         reset.reset_n
		.address       (mm_interconnect_2_timer_1ms_s1_address),    //            s1.address
		.writedata     (mm_interconnect_2_timer_1ms_s1_writedata),  //              .writedata
		.readdata      (mm_interconnect_2_timer_1ms_s1_readdata),   //              .readdata
		.chipselect    (mm_interconnect_2_timer_1ms_s1_chipselect), //              .chipselect
		.write_n       (~mm_interconnect_2_timer_1ms_s1_write),     //              .write_n
		.irq           (irq_synchronizer_receiver_irq),             //           irq.irq
		.timeout_pulse (timer_1ms_external_port_export)             // external_port.export
	);

	MebX_Qsys_Project_timer_1us timer_1us (
		.clk           (clk50_clk),                                 //           clk.clk
		.reset_n       (~rst_controller_019_reset_out_reset),       //         reset.reset_n
		.address       (mm_interconnect_2_timer_1us_s1_address),    //            s1.address
		.writedata     (mm_interconnect_2_timer_1us_s1_writedata),  //              .writedata
		.readdata      (mm_interconnect_2_timer_1us_s1_readdata),   //              .readdata
		.chipselect    (mm_interconnect_2_timer_1us_s1_chipselect), //              .chipselect
		.write_n       (~mm_interconnect_2_timer_1us_s1_write),     //              .write_n
		.irq           (irq_synchronizer_001_receiver_irq),         //           irq.irq
		.timeout_pulse (timer_1us_external_port_export)             // external_port.export
	);

	MebX_Qsys_Project_tristate_conduit_bridge_0 tristate_conduit_bridge_0 (
		.clk                      (m2_ddr2_memory_afi_half_clk_clk),       //   clk.clk
		.reset                    (rst_controller_020_reset_out_reset),    // reset.reset
		.request                  (ext_flash_tcm_request),                 //   tcs.request
		.grant                    (ext_flash_tcm_grant),                   //      .grant
		.tcs_tcm_address_out      (ext_flash_tcm_address_out),             //      .address_out
		.tcs_tcm_read_n_out       (ext_flash_tcm_read_n_out),              //      .read_n_out
		.tcs_tcm_write_n_out      (ext_flash_tcm_write_n_out),             //      .write_n_out
		.tcs_tcm_data_out         (ext_flash_tcm_data_out),                //      .data_out
		.tcs_tcm_data_outen       (ext_flash_tcm_data_outen),              //      .data_outen
		.tcs_tcm_data_in          (ext_flash_tcm_data_in),                 //      .data_in
		.tcs_tcm_chipselect_n_out (ext_flash_tcm_chipselect_n_out),        //      .chipselect_n_out
		.tcm_address_out          (tristate_conduit_tcm_address_out),      //   out.tcm_address_out
		.tcm_read_n_out           (tristate_conduit_tcm_read_n_out),       //      .tcm_read_n_out
		.tcm_write_n_out          (tristate_conduit_tcm_write_n_out),      //      .tcm_write_n_out
		.tcm_data_out             (tristate_conduit_tcm_data_out),         //      .tcm_data_out
		.tcm_chipselect_n_out     (tristate_conduit_tcm_chipselect_n_out)  //      .tcm_chipselect_n_out
	);

	MebX_Qsys_Project_mm_interconnect_0 mm_interconnect_0 (
		.clk_100_clk_clk                                                 (m2_ddr2_memory_afi_half_clk_clk),                                 //                                               clk_100_clk.clk
		.m2_ddr2_memory_afi_clk_clk                                      (m2_ddr2_memory_afi_clk_clk),                                      //                                    m2_ddr2_memory_afi_clk.clk
		.m2_ddr2_memory_afi_half_clk_clk                                 (m2_ddr2_memory_afi_half_clk_clk),                                 //                               m2_ddr2_memory_afi_half_clk.clk
		.COMM_Pedreiro_v1_01_1_reset_sink_reset_bridge_in_reset_reset    (rst_controller_002_reset_out_reset),                              //    COMM_Pedreiro_v1_01_1_reset_sink_reset_bridge_in_reset.reset
		.COMM_Pedreiro_v1_01_2_reset_sink_reset_bridge_in_reset_reset    (rst_controller_003_reset_out_reset),                              //    COMM_Pedreiro_v1_01_2_reset_sink_reset_bridge_in_reset.reset
		.COMM_Pedreiro_v1_01_3_reset_sink_reset_bridge_in_reset_reset    (rst_controller_004_reset_out_reset),                              //    COMM_Pedreiro_v1_01_3_reset_sink_reset_bridge_in_reset.reset
		.COMM_Pedreiro_v1_01_4_reset_sink_reset_bridge_in_reset_reset    (rst_controller_005_reset_out_reset),                              //    COMM_Pedreiro_v1_01_4_reset_sink_reset_bridge_in_reset.reset
		.COMM_Pedreiro_v1_01_5_reset_sink_reset_bridge_in_reset_reset    (rst_controller_006_reset_out_reset),                              //    COMM_Pedreiro_v1_01_5_reset_sink_reset_bridge_in_reset.reset
		.COMM_Pedreiro_v1_01_6_reset_sink_reset_bridge_in_reset_reset    (rst_controller_007_reset_out_reset),                              //    COMM_Pedreiro_v1_01_6_reset_sink_reset_bridge_in_reset.reset
		.FTDI_USB3_0_reset_sink_reset_bridge_in_reset_reset              (rst_controller_008_reset_out_reset),                              //              FTDI_USB3_0_reset_sink_reset_bridge_in_reset.reset
		.m1_clock_bridge_s0_reset_reset_bridge_in_reset_reset            (rst_controller_008_reset_out_reset),                              //            m1_clock_bridge_s0_reset_reset_bridge_in_reset.reset
		.m2_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset (rst_controller_025_reset_out_reset),                              // m2_ddr2_memory_avl_translator_reset_reset_bridge_in_reset.reset
		.m2_ddr2_memory_soft_reset_reset_bridge_in_reset_reset           (rst_controller_025_reset_out_reset),                              //           m2_ddr2_memory_soft_reset_reset_bridge_in_reset.reset
		.COMM_Pedreiro_v1_01_1_avalon_mm_left_buffer_master_address      (comm_pedreiro_v1_01_1_avalon_mm_left_buffer_master_address),      //        COMM_Pedreiro_v1_01_1_avalon_mm_left_buffer_master.address
		.COMM_Pedreiro_v1_01_1_avalon_mm_left_buffer_master_waitrequest  (comm_pedreiro_v1_01_1_avalon_mm_left_buffer_master_waitrequest),  //                                                          .waitrequest
		.COMM_Pedreiro_v1_01_1_avalon_mm_left_buffer_master_read         (comm_pedreiro_v1_01_1_avalon_mm_left_buffer_master_read),         //                                                          .read
		.COMM_Pedreiro_v1_01_1_avalon_mm_left_buffer_master_readdata     (comm_pedreiro_v1_01_1_avalon_mm_left_buffer_master_readdata),     //                                                          .readdata
		.COMM_Pedreiro_v1_01_1_avalon_mm_right_buffer_master_address     (comm_pedreiro_v1_01_1_avalon_mm_right_buffer_master_address),     //       COMM_Pedreiro_v1_01_1_avalon_mm_right_buffer_master.address
		.COMM_Pedreiro_v1_01_1_avalon_mm_right_buffer_master_waitrequest (comm_pedreiro_v1_01_1_avalon_mm_right_buffer_master_waitrequest), //                                                          .waitrequest
		.COMM_Pedreiro_v1_01_1_avalon_mm_right_buffer_master_read        (comm_pedreiro_v1_01_1_avalon_mm_right_buffer_master_read),        //                                                          .read
		.COMM_Pedreiro_v1_01_1_avalon_mm_right_buffer_master_readdata    (comm_pedreiro_v1_01_1_avalon_mm_right_buffer_master_readdata),    //                                                          .readdata
		.COMM_Pedreiro_v1_01_2_avalon_mm_left_buffer_master_address      (comm_pedreiro_v1_01_2_avalon_mm_left_buffer_master_address),      //        COMM_Pedreiro_v1_01_2_avalon_mm_left_buffer_master.address
		.COMM_Pedreiro_v1_01_2_avalon_mm_left_buffer_master_waitrequest  (comm_pedreiro_v1_01_2_avalon_mm_left_buffer_master_waitrequest),  //                                                          .waitrequest
		.COMM_Pedreiro_v1_01_2_avalon_mm_left_buffer_master_read         (comm_pedreiro_v1_01_2_avalon_mm_left_buffer_master_read),         //                                                          .read
		.COMM_Pedreiro_v1_01_2_avalon_mm_left_buffer_master_readdata     (comm_pedreiro_v1_01_2_avalon_mm_left_buffer_master_readdata),     //                                                          .readdata
		.COMM_Pedreiro_v1_01_2_avalon_mm_right_buffer_master_address     (comm_pedreiro_v1_01_2_avalon_mm_right_buffer_master_address),     //       COMM_Pedreiro_v1_01_2_avalon_mm_right_buffer_master.address
		.COMM_Pedreiro_v1_01_2_avalon_mm_right_buffer_master_waitrequest (comm_pedreiro_v1_01_2_avalon_mm_right_buffer_master_waitrequest), //                                                          .waitrequest
		.COMM_Pedreiro_v1_01_2_avalon_mm_right_buffer_master_read        (comm_pedreiro_v1_01_2_avalon_mm_right_buffer_master_read),        //                                                          .read
		.COMM_Pedreiro_v1_01_2_avalon_mm_right_buffer_master_readdata    (comm_pedreiro_v1_01_2_avalon_mm_right_buffer_master_readdata),    //                                                          .readdata
		.COMM_Pedreiro_v1_01_3_avalon_mm_left_buffer_master_address      (comm_pedreiro_v1_01_3_avalon_mm_left_buffer_master_address),      //        COMM_Pedreiro_v1_01_3_avalon_mm_left_buffer_master.address
		.COMM_Pedreiro_v1_01_3_avalon_mm_left_buffer_master_waitrequest  (comm_pedreiro_v1_01_3_avalon_mm_left_buffer_master_waitrequest),  //                                                          .waitrequest
		.COMM_Pedreiro_v1_01_3_avalon_mm_left_buffer_master_read         (comm_pedreiro_v1_01_3_avalon_mm_left_buffer_master_read),         //                                                          .read
		.COMM_Pedreiro_v1_01_3_avalon_mm_left_buffer_master_readdata     (comm_pedreiro_v1_01_3_avalon_mm_left_buffer_master_readdata),     //                                                          .readdata
		.COMM_Pedreiro_v1_01_3_avalon_mm_right_buffer_master_address     (comm_pedreiro_v1_01_3_avalon_mm_right_buffer_master_address),     //       COMM_Pedreiro_v1_01_3_avalon_mm_right_buffer_master.address
		.COMM_Pedreiro_v1_01_3_avalon_mm_right_buffer_master_waitrequest (comm_pedreiro_v1_01_3_avalon_mm_right_buffer_master_waitrequest), //                                                          .waitrequest
		.COMM_Pedreiro_v1_01_3_avalon_mm_right_buffer_master_read        (comm_pedreiro_v1_01_3_avalon_mm_right_buffer_master_read),        //                                                          .read
		.COMM_Pedreiro_v1_01_3_avalon_mm_right_buffer_master_readdata    (comm_pedreiro_v1_01_3_avalon_mm_right_buffer_master_readdata),    //                                                          .readdata
		.COMM_Pedreiro_v1_01_4_avalon_mm_left_buffer_master_address      (comm_pedreiro_v1_01_4_avalon_mm_left_buffer_master_address),      //        COMM_Pedreiro_v1_01_4_avalon_mm_left_buffer_master.address
		.COMM_Pedreiro_v1_01_4_avalon_mm_left_buffer_master_waitrequest  (comm_pedreiro_v1_01_4_avalon_mm_left_buffer_master_waitrequest),  //                                                          .waitrequest
		.COMM_Pedreiro_v1_01_4_avalon_mm_left_buffer_master_read         (comm_pedreiro_v1_01_4_avalon_mm_left_buffer_master_read),         //                                                          .read
		.COMM_Pedreiro_v1_01_4_avalon_mm_left_buffer_master_readdata     (comm_pedreiro_v1_01_4_avalon_mm_left_buffer_master_readdata),     //                                                          .readdata
		.COMM_Pedreiro_v1_01_4_avalon_mm_right_buffer_master_address     (comm_pedreiro_v1_01_4_avalon_mm_right_buffer_master_address),     //       COMM_Pedreiro_v1_01_4_avalon_mm_right_buffer_master.address
		.COMM_Pedreiro_v1_01_4_avalon_mm_right_buffer_master_waitrequest (comm_pedreiro_v1_01_4_avalon_mm_right_buffer_master_waitrequest), //                                                          .waitrequest
		.COMM_Pedreiro_v1_01_4_avalon_mm_right_buffer_master_read        (comm_pedreiro_v1_01_4_avalon_mm_right_buffer_master_read),        //                                                          .read
		.COMM_Pedreiro_v1_01_4_avalon_mm_right_buffer_master_readdata    (comm_pedreiro_v1_01_4_avalon_mm_right_buffer_master_readdata),    //                                                          .readdata
		.COMM_Pedreiro_v1_01_5_avalon_mm_left_buffer_master_address      (comm_pedreiro_v1_01_5_avalon_mm_left_buffer_master_address),      //        COMM_Pedreiro_v1_01_5_avalon_mm_left_buffer_master.address
		.COMM_Pedreiro_v1_01_5_avalon_mm_left_buffer_master_waitrequest  (comm_pedreiro_v1_01_5_avalon_mm_left_buffer_master_waitrequest),  //                                                          .waitrequest
		.COMM_Pedreiro_v1_01_5_avalon_mm_left_buffer_master_read         (comm_pedreiro_v1_01_5_avalon_mm_left_buffer_master_read),         //                                                          .read
		.COMM_Pedreiro_v1_01_5_avalon_mm_left_buffer_master_readdata     (comm_pedreiro_v1_01_5_avalon_mm_left_buffer_master_readdata),     //                                                          .readdata
		.COMM_Pedreiro_v1_01_5_avalon_mm_right_buffer_master_address     (comm_pedreiro_v1_01_5_avalon_mm_right_buffer_master_address),     //       COMM_Pedreiro_v1_01_5_avalon_mm_right_buffer_master.address
		.COMM_Pedreiro_v1_01_5_avalon_mm_right_buffer_master_waitrequest (comm_pedreiro_v1_01_5_avalon_mm_right_buffer_master_waitrequest), //                                                          .waitrequest
		.COMM_Pedreiro_v1_01_5_avalon_mm_right_buffer_master_read        (comm_pedreiro_v1_01_5_avalon_mm_right_buffer_master_read),        //                                                          .read
		.COMM_Pedreiro_v1_01_5_avalon_mm_right_buffer_master_readdata    (comm_pedreiro_v1_01_5_avalon_mm_right_buffer_master_readdata),    //                                                          .readdata
		.COMM_Pedreiro_v1_01_6_avalon_mm_left_buffer_master_address      (comm_pedreiro_v1_01_6_avalon_mm_left_buffer_master_address),      //        COMM_Pedreiro_v1_01_6_avalon_mm_left_buffer_master.address
		.COMM_Pedreiro_v1_01_6_avalon_mm_left_buffer_master_waitrequest  (comm_pedreiro_v1_01_6_avalon_mm_left_buffer_master_waitrequest),  //                                                          .waitrequest
		.COMM_Pedreiro_v1_01_6_avalon_mm_left_buffer_master_read         (comm_pedreiro_v1_01_6_avalon_mm_left_buffer_master_read),         //                                                          .read
		.COMM_Pedreiro_v1_01_6_avalon_mm_left_buffer_master_readdata     (comm_pedreiro_v1_01_6_avalon_mm_left_buffer_master_readdata),     //                                                          .readdata
		.COMM_Pedreiro_v1_01_6_avalon_mm_right_buffer_master_address     (comm_pedreiro_v1_01_6_avalon_mm_right_buffer_master_address),     //       COMM_Pedreiro_v1_01_6_avalon_mm_right_buffer_master.address
		.COMM_Pedreiro_v1_01_6_avalon_mm_right_buffer_master_waitrequest (comm_pedreiro_v1_01_6_avalon_mm_right_buffer_master_waitrequest), //                                                          .waitrequest
		.COMM_Pedreiro_v1_01_6_avalon_mm_right_buffer_master_read        (comm_pedreiro_v1_01_6_avalon_mm_right_buffer_master_read),        //                                                          .read
		.COMM_Pedreiro_v1_01_6_avalon_mm_right_buffer_master_readdata    (comm_pedreiro_v1_01_6_avalon_mm_right_buffer_master_readdata),    //                                                          .readdata
		.ddr2_address_span_extender_expanded_master_address              (ddr2_address_span_extender_expanded_master_address),              //                ddr2_address_span_extender_expanded_master.address
		.ddr2_address_span_extender_expanded_master_waitrequest          (ddr2_address_span_extender_expanded_master_waitrequest),          //                                                          .waitrequest
		.ddr2_address_span_extender_expanded_master_burstcount           (ddr2_address_span_extender_expanded_master_burstcount),           //                                                          .burstcount
		.ddr2_address_span_extender_expanded_master_byteenable           (ddr2_address_span_extender_expanded_master_byteenable),           //                                                          .byteenable
		.ddr2_address_span_extender_expanded_master_read                 (ddr2_address_span_extender_expanded_master_read),                 //                                                          .read
		.ddr2_address_span_extender_expanded_master_readdata             (ddr2_address_span_extender_expanded_master_readdata),             //                                                          .readdata
		.ddr2_address_span_extender_expanded_master_readdatavalid        (ddr2_address_span_extender_expanded_master_readdatavalid),        //                                                          .readdatavalid
		.ddr2_address_span_extender_expanded_master_write                (ddr2_address_span_extender_expanded_master_write),                //                                                          .write
		.ddr2_address_span_extender_expanded_master_writedata            (ddr2_address_span_extender_expanded_master_writedata),            //                                                          .writedata
		.FTDI_USB3_0_avalon_master_data_address                          (ftdi_usb3_0_avalon_master_data_address),                          //                            FTDI_USB3_0_avalon_master_data.address
		.FTDI_USB3_0_avalon_master_data_waitrequest                      (ftdi_usb3_0_avalon_master_data_waitrequest),                      //                                                          .waitrequest
		.FTDI_USB3_0_avalon_master_data_read                             (ftdi_usb3_0_avalon_master_data_read),                             //                                                          .read
		.FTDI_USB3_0_avalon_master_data_readdata                         (ftdi_usb3_0_avalon_master_data_readdata),                         //                                                          .readdata
		.FTDI_USB3_0_avalon_master_data_write                            (ftdi_usb3_0_avalon_master_data_write),                            //                                                          .write
		.FTDI_USB3_0_avalon_master_data_writedata                        (ftdi_usb3_0_avalon_master_data_writedata),                        //                                                          .writedata
		.rmap_mem_nfee_comm_1_avalon_mm_rmap_master_address              (rmap_mem_nfee_comm_1_avalon_mm_rmap_master_address),              //                rmap_mem_nfee_comm_1_avalon_mm_rmap_master.address
		.rmap_mem_nfee_comm_1_avalon_mm_rmap_master_waitrequest          (rmap_mem_nfee_comm_1_avalon_mm_rmap_master_waitrequest),          //                                                          .waitrequest
		.rmap_mem_nfee_comm_1_avalon_mm_rmap_master_read                 (rmap_mem_nfee_comm_1_avalon_mm_rmap_master_read),                 //                                                          .read
		.rmap_mem_nfee_comm_1_avalon_mm_rmap_master_readdata             (rmap_mem_nfee_comm_1_avalon_mm_rmap_master_readdata),             //                                                          .readdata
		.rmap_mem_nfee_comm_1_avalon_mm_rmap_master_write                (rmap_mem_nfee_comm_1_avalon_mm_rmap_master_write),                //                                                          .write
		.rmap_mem_nfee_comm_1_avalon_mm_rmap_master_writedata            (rmap_mem_nfee_comm_1_avalon_mm_rmap_master_writedata),            //                                                          .writedata
		.rmap_mem_nfee_comm_2_avalon_mm_rmap_master_address              (rmap_mem_nfee_comm_2_avalon_mm_rmap_master_address),              //                rmap_mem_nfee_comm_2_avalon_mm_rmap_master.address
		.rmap_mem_nfee_comm_2_avalon_mm_rmap_master_waitrequest          (rmap_mem_nfee_comm_2_avalon_mm_rmap_master_waitrequest),          //                                                          .waitrequest
		.rmap_mem_nfee_comm_2_avalon_mm_rmap_master_read                 (rmap_mem_nfee_comm_2_avalon_mm_rmap_master_read),                 //                                                          .read
		.rmap_mem_nfee_comm_2_avalon_mm_rmap_master_readdata             (rmap_mem_nfee_comm_2_avalon_mm_rmap_master_readdata),             //                                                          .readdata
		.rmap_mem_nfee_comm_2_avalon_mm_rmap_master_write                (rmap_mem_nfee_comm_2_avalon_mm_rmap_master_write),                //                                                          .write
		.rmap_mem_nfee_comm_2_avalon_mm_rmap_master_writedata            (rmap_mem_nfee_comm_2_avalon_mm_rmap_master_writedata),            //                                                          .writedata
		.rmap_mem_nfee_comm_3_avalon_mm_rmap_master_address              (rmap_mem_nfee_comm_3_avalon_mm_rmap_master_address),              //                rmap_mem_nfee_comm_3_avalon_mm_rmap_master.address
		.rmap_mem_nfee_comm_3_avalon_mm_rmap_master_waitrequest          (rmap_mem_nfee_comm_3_avalon_mm_rmap_master_waitrequest),          //                                                          .waitrequest
		.rmap_mem_nfee_comm_3_avalon_mm_rmap_master_read                 (rmap_mem_nfee_comm_3_avalon_mm_rmap_master_read),                 //                                                          .read
		.rmap_mem_nfee_comm_3_avalon_mm_rmap_master_readdata             (rmap_mem_nfee_comm_3_avalon_mm_rmap_master_readdata),             //                                                          .readdata
		.rmap_mem_nfee_comm_3_avalon_mm_rmap_master_write                (rmap_mem_nfee_comm_3_avalon_mm_rmap_master_write),                //                                                          .write
		.rmap_mem_nfee_comm_3_avalon_mm_rmap_master_writedata            (rmap_mem_nfee_comm_3_avalon_mm_rmap_master_writedata),            //                                                          .writedata
		.rmap_mem_nfee_comm_4_avalon_mm_rmap_master_address              (rmap_mem_nfee_comm_4_avalon_mm_rmap_master_address),              //                rmap_mem_nfee_comm_4_avalon_mm_rmap_master.address
		.rmap_mem_nfee_comm_4_avalon_mm_rmap_master_waitrequest          (rmap_mem_nfee_comm_4_avalon_mm_rmap_master_waitrequest),          //                                                          .waitrequest
		.rmap_mem_nfee_comm_4_avalon_mm_rmap_master_read                 (rmap_mem_nfee_comm_4_avalon_mm_rmap_master_read),                 //                                                          .read
		.rmap_mem_nfee_comm_4_avalon_mm_rmap_master_readdata             (rmap_mem_nfee_comm_4_avalon_mm_rmap_master_readdata),             //                                                          .readdata
		.rmap_mem_nfee_comm_4_avalon_mm_rmap_master_write                (rmap_mem_nfee_comm_4_avalon_mm_rmap_master_write),                //                                                          .write
		.rmap_mem_nfee_comm_4_avalon_mm_rmap_master_writedata            (rmap_mem_nfee_comm_4_avalon_mm_rmap_master_writedata),            //                                                          .writedata
		.rmap_mem_nfee_comm_5_avalon_mm_rmap_master_address              (rmap_mem_nfee_comm_5_avalon_mm_rmap_master_address),              //                rmap_mem_nfee_comm_5_avalon_mm_rmap_master.address
		.rmap_mem_nfee_comm_5_avalon_mm_rmap_master_waitrequest          (rmap_mem_nfee_comm_5_avalon_mm_rmap_master_waitrequest),          //                                                          .waitrequest
		.rmap_mem_nfee_comm_5_avalon_mm_rmap_master_read                 (rmap_mem_nfee_comm_5_avalon_mm_rmap_master_read),                 //                                                          .read
		.rmap_mem_nfee_comm_5_avalon_mm_rmap_master_readdata             (rmap_mem_nfee_comm_5_avalon_mm_rmap_master_readdata),             //                                                          .readdata
		.rmap_mem_nfee_comm_5_avalon_mm_rmap_master_write                (rmap_mem_nfee_comm_5_avalon_mm_rmap_master_write),                //                                                          .write
		.rmap_mem_nfee_comm_5_avalon_mm_rmap_master_writedata            (rmap_mem_nfee_comm_5_avalon_mm_rmap_master_writedata),            //                                                          .writedata
		.rmap_mem_nfee_comm_6_avalon_mm_rmap_master_address              (rmap_mem_nfee_comm_6_avalon_mm_rmap_master_address),              //                rmap_mem_nfee_comm_6_avalon_mm_rmap_master.address
		.rmap_mem_nfee_comm_6_avalon_mm_rmap_master_waitrequest          (rmap_mem_nfee_comm_6_avalon_mm_rmap_master_waitrequest),          //                                                          .waitrequest
		.rmap_mem_nfee_comm_6_avalon_mm_rmap_master_read                 (rmap_mem_nfee_comm_6_avalon_mm_rmap_master_read),                 //                                                          .read
		.rmap_mem_nfee_comm_6_avalon_mm_rmap_master_readdata             (rmap_mem_nfee_comm_6_avalon_mm_rmap_master_readdata),             //                                                          .readdata
		.rmap_mem_nfee_comm_6_avalon_mm_rmap_master_write                (rmap_mem_nfee_comm_6_avalon_mm_rmap_master_write),                //                                                          .write
		.rmap_mem_nfee_comm_6_avalon_mm_rmap_master_writedata            (rmap_mem_nfee_comm_6_avalon_mm_rmap_master_writedata),            //                                                          .writedata
		.m1_clock_bridge_s0_address                                      (mm_interconnect_0_m1_clock_bridge_s0_address),                    //                                        m1_clock_bridge_s0.address
		.m1_clock_bridge_s0_write                                        (mm_interconnect_0_m1_clock_bridge_s0_write),                      //                                                          .write
		.m1_clock_bridge_s0_read                                         (mm_interconnect_0_m1_clock_bridge_s0_read),                       //                                                          .read
		.m1_clock_bridge_s0_readdata                                     (mm_interconnect_0_m1_clock_bridge_s0_readdata),                   //                                                          .readdata
		.m1_clock_bridge_s0_writedata                                    (mm_interconnect_0_m1_clock_bridge_s0_writedata),                  //                                                          .writedata
		.m1_clock_bridge_s0_burstcount                                   (mm_interconnect_0_m1_clock_bridge_s0_burstcount),                 //                                                          .burstcount
		.m1_clock_bridge_s0_byteenable                                   (mm_interconnect_0_m1_clock_bridge_s0_byteenable),                 //                                                          .byteenable
		.m1_clock_bridge_s0_readdatavalid                                (mm_interconnect_0_m1_clock_bridge_s0_readdatavalid),              //                                                          .readdatavalid
		.m1_clock_bridge_s0_waitrequest                                  (mm_interconnect_0_m1_clock_bridge_s0_waitrequest),                //                                                          .waitrequest
		.m1_clock_bridge_s0_debugaccess                                  (mm_interconnect_0_m1_clock_bridge_s0_debugaccess),                //                                                          .debugaccess
		.m2_ddr2_memory_avl_address                                      (mm_interconnect_0_m2_ddr2_memory_avl_address),                    //                                        m2_ddr2_memory_avl.address
		.m2_ddr2_memory_avl_write                                        (mm_interconnect_0_m2_ddr2_memory_avl_write),                      //                                                          .write
		.m2_ddr2_memory_avl_read                                         (mm_interconnect_0_m2_ddr2_memory_avl_read),                       //                                                          .read
		.m2_ddr2_memory_avl_readdata                                     (mm_interconnect_0_m2_ddr2_memory_avl_readdata),                   //                                                          .readdata
		.m2_ddr2_memory_avl_writedata                                    (mm_interconnect_0_m2_ddr2_memory_avl_writedata),                  //                                                          .writedata
		.m2_ddr2_memory_avl_beginbursttransfer                           (mm_interconnect_0_m2_ddr2_memory_avl_beginbursttransfer),         //                                                          .beginbursttransfer
		.m2_ddr2_memory_avl_burstcount                                   (mm_interconnect_0_m2_ddr2_memory_avl_burstcount),                 //                                                          .burstcount
		.m2_ddr2_memory_avl_byteenable                                   (mm_interconnect_0_m2_ddr2_memory_avl_byteenable),                 //                                                          .byteenable
		.m2_ddr2_memory_avl_readdatavalid                                (mm_interconnect_0_m2_ddr2_memory_avl_readdatavalid),              //                                                          .readdatavalid
		.m2_ddr2_memory_avl_waitrequest                                  (~mm_interconnect_0_m2_ddr2_memory_avl_waitrequest)                //                                                          .waitrequest
	);

	MebX_Qsys_Project_mm_interconnect_1 mm_interconnect_1 (
		.clk_100_clk_clk                                             (m2_ddr2_memory_afi_half_clk_clk),                                            //                                           clk_100_clk.clk
		.ext_flash_reset_reset_bridge_in_reset_reset                 (rst_controller_020_reset_out_reset),                                         //                 ext_flash_reset_reset_bridge_in_reset.reset
		.jtag_uart_0_reset_reset_bridge_in_reset_reset               (rst_controller_008_reset_out_reset),                                         //               jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset              (rst_controller_022_reset_out_reset),                                         //              nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.rmap_mem_nfee_comm_1_reset_sink_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                         // rmap_mem_nfee_comm_1_reset_sink_reset_bridge_in_reset.reset
		.rmap_mem_nfee_comm_2_reset_sink_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                                         // rmap_mem_nfee_comm_2_reset_sink_reset_bridge_in_reset.reset
		.rmap_mem_nfee_comm_3_reset_sink_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                                         // rmap_mem_nfee_comm_3_reset_sink_reset_bridge_in_reset.reset
		.rmap_mem_nfee_comm_4_reset_sink_reset_bridge_in_reset_reset (rst_controller_005_reset_out_reset),                                         // rmap_mem_nfee_comm_4_reset_sink_reset_bridge_in_reset.reset
		.rmap_mem_nfee_comm_5_reset_sink_reset_bridge_in_reset_reset (rst_controller_006_reset_out_reset),                                         // rmap_mem_nfee_comm_5_reset_sink_reset_bridge_in_reset.reset
		.rmap_mem_nfee_comm_6_reset_sink_reset_bridge_in_reset_reset (rst_controller_007_reset_out_reset),                                         // rmap_mem_nfee_comm_6_reset_sink_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                            (nios2_gen2_0_data_master_address),                                           //                              nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                        (nios2_gen2_0_data_master_waitrequest),                                       //                                                      .waitrequest
		.nios2_gen2_0_data_master_byteenable                         (nios2_gen2_0_data_master_byteenable),                                        //                                                      .byteenable
		.nios2_gen2_0_data_master_read                               (nios2_gen2_0_data_master_read),                                              //                                                      .read
		.nios2_gen2_0_data_master_readdata                           (nios2_gen2_0_data_master_readdata),                                          //                                                      .readdata
		.nios2_gen2_0_data_master_write                              (nios2_gen2_0_data_master_write),                                             //                                                      .write
		.nios2_gen2_0_data_master_writedata                          (nios2_gen2_0_data_master_writedata),                                         //                                                      .writedata
		.nios2_gen2_0_data_master_debugaccess                        (nios2_gen2_0_data_master_debugaccess),                                       //                                                      .debugaccess
		.nios2_gen2_0_instruction_master_address                     (nios2_gen2_0_instruction_master_address),                                    //                       nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                 (nios2_gen2_0_instruction_master_waitrequest),                                //                                                      .waitrequest
		.nios2_gen2_0_instruction_master_burstcount                  (nios2_gen2_0_instruction_master_burstcount),                                 //                                                      .burstcount
		.nios2_gen2_0_instruction_master_read                        (nios2_gen2_0_instruction_master_read),                                       //                                                      .read
		.nios2_gen2_0_instruction_master_readdata                    (nios2_gen2_0_instruction_master_readdata),                                   //                                                      .readdata
		.nios2_gen2_0_instruction_master_readdatavalid               (nios2_gen2_0_instruction_master_readdatavalid),                              //                                                      .readdatavalid
		.clock_bridge_afi_50_s0_address                              (mm_interconnect_1_clock_bridge_afi_50_s0_address),                           //                                clock_bridge_afi_50_s0.address
		.clock_bridge_afi_50_s0_write                                (mm_interconnect_1_clock_bridge_afi_50_s0_write),                             //                                                      .write
		.clock_bridge_afi_50_s0_read                                 (mm_interconnect_1_clock_bridge_afi_50_s0_read),                              //                                                      .read
		.clock_bridge_afi_50_s0_readdata                             (mm_interconnect_1_clock_bridge_afi_50_s0_readdata),                          //                                                      .readdata
		.clock_bridge_afi_50_s0_writedata                            (mm_interconnect_1_clock_bridge_afi_50_s0_writedata),                         //                                                      .writedata
		.clock_bridge_afi_50_s0_burstcount                           (mm_interconnect_1_clock_bridge_afi_50_s0_burstcount),                        //                                                      .burstcount
		.clock_bridge_afi_50_s0_byteenable                           (mm_interconnect_1_clock_bridge_afi_50_s0_byteenable),                        //                                                      .byteenable
		.clock_bridge_afi_50_s0_readdatavalid                        (mm_interconnect_1_clock_bridge_afi_50_s0_readdatavalid),                     //                                                      .readdatavalid
		.clock_bridge_afi_50_s0_waitrequest                          (mm_interconnect_1_clock_bridge_afi_50_s0_waitrequest),                       //                                                      .waitrequest
		.clock_bridge_afi_50_s0_debugaccess                          (mm_interconnect_1_clock_bridge_afi_50_s0_debugaccess),                       //                                                      .debugaccess
		.COMM_Pedreiro_v1_01_1_avalon_slave_windowing_address        (mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_address),     //          COMM_Pedreiro_v1_01_1_avalon_slave_windowing.address
		.COMM_Pedreiro_v1_01_1_avalon_slave_windowing_write          (mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_write),       //                                                      .write
		.COMM_Pedreiro_v1_01_1_avalon_slave_windowing_read           (mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_read),        //                                                      .read
		.COMM_Pedreiro_v1_01_1_avalon_slave_windowing_readdata       (mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_readdata),    //                                                      .readdata
		.COMM_Pedreiro_v1_01_1_avalon_slave_windowing_writedata      (mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_writedata),   //                                                      .writedata
		.COMM_Pedreiro_v1_01_1_avalon_slave_windowing_byteenable     (mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_byteenable),  //                                                      .byteenable
		.COMM_Pedreiro_v1_01_1_avalon_slave_windowing_waitrequest    (mm_interconnect_1_comm_pedreiro_v1_01_1_avalon_slave_windowing_waitrequest), //                                                      .waitrequest
		.COMM_Pedreiro_v1_01_2_avalon_slave_windowing_address        (mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_address),     //          COMM_Pedreiro_v1_01_2_avalon_slave_windowing.address
		.COMM_Pedreiro_v1_01_2_avalon_slave_windowing_write          (mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_write),       //                                                      .write
		.COMM_Pedreiro_v1_01_2_avalon_slave_windowing_read           (mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_read),        //                                                      .read
		.COMM_Pedreiro_v1_01_2_avalon_slave_windowing_readdata       (mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_readdata),    //                                                      .readdata
		.COMM_Pedreiro_v1_01_2_avalon_slave_windowing_writedata      (mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_writedata),   //                                                      .writedata
		.COMM_Pedreiro_v1_01_2_avalon_slave_windowing_byteenable     (mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_byteenable),  //                                                      .byteenable
		.COMM_Pedreiro_v1_01_2_avalon_slave_windowing_waitrequest    (mm_interconnect_1_comm_pedreiro_v1_01_2_avalon_slave_windowing_waitrequest), //                                                      .waitrequest
		.COMM_Pedreiro_v1_01_3_avalon_slave_windowing_address        (mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_address),     //          COMM_Pedreiro_v1_01_3_avalon_slave_windowing.address
		.COMM_Pedreiro_v1_01_3_avalon_slave_windowing_write          (mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_write),       //                                                      .write
		.COMM_Pedreiro_v1_01_3_avalon_slave_windowing_read           (mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_read),        //                                                      .read
		.COMM_Pedreiro_v1_01_3_avalon_slave_windowing_readdata       (mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_readdata),    //                                                      .readdata
		.COMM_Pedreiro_v1_01_3_avalon_slave_windowing_writedata      (mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_writedata),   //                                                      .writedata
		.COMM_Pedreiro_v1_01_3_avalon_slave_windowing_byteenable     (mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_byteenable),  //                                                      .byteenable
		.COMM_Pedreiro_v1_01_3_avalon_slave_windowing_waitrequest    (mm_interconnect_1_comm_pedreiro_v1_01_3_avalon_slave_windowing_waitrequest), //                                                      .waitrequest
		.COMM_Pedreiro_v1_01_4_avalon_slave_windowing_address        (mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_address),     //          COMM_Pedreiro_v1_01_4_avalon_slave_windowing.address
		.COMM_Pedreiro_v1_01_4_avalon_slave_windowing_write          (mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_write),       //                                                      .write
		.COMM_Pedreiro_v1_01_4_avalon_slave_windowing_read           (mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_read),        //                                                      .read
		.COMM_Pedreiro_v1_01_4_avalon_slave_windowing_readdata       (mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_readdata),    //                                                      .readdata
		.COMM_Pedreiro_v1_01_4_avalon_slave_windowing_writedata      (mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_writedata),   //                                                      .writedata
		.COMM_Pedreiro_v1_01_4_avalon_slave_windowing_byteenable     (mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_byteenable),  //                                                      .byteenable
		.COMM_Pedreiro_v1_01_4_avalon_slave_windowing_waitrequest    (mm_interconnect_1_comm_pedreiro_v1_01_4_avalon_slave_windowing_waitrequest), //                                                      .waitrequest
		.COMM_Pedreiro_v1_01_5_avalon_slave_windowing_address        (mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_address),     //          COMM_Pedreiro_v1_01_5_avalon_slave_windowing.address
		.COMM_Pedreiro_v1_01_5_avalon_slave_windowing_write          (mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_write),       //                                                      .write
		.COMM_Pedreiro_v1_01_5_avalon_slave_windowing_read           (mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_read),        //                                                      .read
		.COMM_Pedreiro_v1_01_5_avalon_slave_windowing_readdata       (mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_readdata),    //                                                      .readdata
		.COMM_Pedreiro_v1_01_5_avalon_slave_windowing_writedata      (mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_writedata),   //                                                      .writedata
		.COMM_Pedreiro_v1_01_5_avalon_slave_windowing_byteenable     (mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_byteenable),  //                                                      .byteenable
		.COMM_Pedreiro_v1_01_5_avalon_slave_windowing_waitrequest    (mm_interconnect_1_comm_pedreiro_v1_01_5_avalon_slave_windowing_waitrequest), //                                                      .waitrequest
		.COMM_Pedreiro_v1_01_6_avalon_slave_windowing_address        (mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_address),     //          COMM_Pedreiro_v1_01_6_avalon_slave_windowing.address
		.COMM_Pedreiro_v1_01_6_avalon_slave_windowing_write          (mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_write),       //                                                      .write
		.COMM_Pedreiro_v1_01_6_avalon_slave_windowing_read           (mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_read),        //                                                      .read
		.COMM_Pedreiro_v1_01_6_avalon_slave_windowing_readdata       (mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_readdata),    //                                                      .readdata
		.COMM_Pedreiro_v1_01_6_avalon_slave_windowing_writedata      (mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_writedata),   //                                                      .writedata
		.COMM_Pedreiro_v1_01_6_avalon_slave_windowing_byteenable     (mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_byteenable),  //                                                      .byteenable
		.COMM_Pedreiro_v1_01_6_avalon_slave_windowing_waitrequest    (mm_interconnect_1_comm_pedreiro_v1_01_6_avalon_slave_windowing_waitrequest), //                                                      .waitrequest
		.ddr2_address_span_extender_cntl_write                       (mm_interconnect_1_ddr2_address_span_extender_cntl_write),                    //                       ddr2_address_span_extender_cntl.write
		.ddr2_address_span_extender_cntl_read                        (mm_interconnect_1_ddr2_address_span_extender_cntl_read),                     //                                                      .read
		.ddr2_address_span_extender_cntl_readdata                    (mm_interconnect_1_ddr2_address_span_extender_cntl_readdata),                 //                                                      .readdata
		.ddr2_address_span_extender_cntl_writedata                   (mm_interconnect_1_ddr2_address_span_extender_cntl_writedata),                //                                                      .writedata
		.ddr2_address_span_extender_cntl_byteenable                  (mm_interconnect_1_ddr2_address_span_extender_cntl_byteenable),               //                                                      .byteenable
		.ddr2_address_span_extender_windowed_slave_address           (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_address),        //             ddr2_address_span_extender_windowed_slave.address
		.ddr2_address_span_extender_windowed_slave_write             (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_write),          //                                                      .write
		.ddr2_address_span_extender_windowed_slave_read              (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_read),           //                                                      .read
		.ddr2_address_span_extender_windowed_slave_readdata          (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdata),       //                                                      .readdata
		.ddr2_address_span_extender_windowed_slave_writedata         (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_writedata),      //                                                      .writedata
		.ddr2_address_span_extender_windowed_slave_burstcount        (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_burstcount),     //                                                      .burstcount
		.ddr2_address_span_extender_windowed_slave_byteenable        (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_byteenable),     //                                                      .byteenable
		.ddr2_address_span_extender_windowed_slave_readdatavalid     (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdatavalid),  //                                                      .readdatavalid
		.ddr2_address_span_extender_windowed_slave_waitrequest       (mm_interconnect_1_ddr2_address_span_extender_windowed_slave_waitrequest),    //                                                      .waitrequest
		.ext_flash_uas_address                                       (mm_interconnect_1_ext_flash_uas_address),                                    //                                         ext_flash_uas.address
		.ext_flash_uas_write                                         (mm_interconnect_1_ext_flash_uas_write),                                      //                                                      .write
		.ext_flash_uas_read                                          (mm_interconnect_1_ext_flash_uas_read),                                       //                                                      .read
		.ext_flash_uas_readdata                                      (mm_interconnect_1_ext_flash_uas_readdata),                                   //                                                      .readdata
		.ext_flash_uas_writedata                                     (mm_interconnect_1_ext_flash_uas_writedata),                                  //                                                      .writedata
		.ext_flash_uas_burstcount                                    (mm_interconnect_1_ext_flash_uas_burstcount),                                 //                                                      .burstcount
		.ext_flash_uas_byteenable                                    (mm_interconnect_1_ext_flash_uas_byteenable),                                 //                                                      .byteenable
		.ext_flash_uas_readdatavalid                                 (mm_interconnect_1_ext_flash_uas_readdatavalid),                              //                                                      .readdatavalid
		.ext_flash_uas_waitrequest                                   (mm_interconnect_1_ext_flash_uas_waitrequest),                                //                                                      .waitrequest
		.ext_flash_uas_lock                                          (mm_interconnect_1_ext_flash_uas_lock),                                       //                                                      .lock
		.ext_flash_uas_debugaccess                                   (mm_interconnect_1_ext_flash_uas_debugaccess),                                //                                                      .debugaccess
		.FTDI_USB3_0_avalon_slave_config_address                     (mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_address),                  //                       FTDI_USB3_0_avalon_slave_config.address
		.FTDI_USB3_0_avalon_slave_config_write                       (mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_write),                    //                                                      .write
		.FTDI_USB3_0_avalon_slave_config_read                        (mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_read),                     //                                                      .read
		.FTDI_USB3_0_avalon_slave_config_readdata                    (mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_readdata),                 //                                                      .readdata
		.FTDI_USB3_0_avalon_slave_config_writedata                   (mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_writedata),                //                                                      .writedata
		.FTDI_USB3_0_avalon_slave_config_byteenable                  (mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_byteenable),               //                                                      .byteenable
		.FTDI_USB3_0_avalon_slave_config_waitrequest                 (mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_waitrequest),              //                                                      .waitrequest
		.jtag_uart_0_avalon_jtag_slave_address                       (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),                    //                         jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                         (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),                      //                                                      .write
		.jtag_uart_0_avalon_jtag_slave_read                          (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),                       //                                                      .read
		.jtag_uart_0_avalon_jtag_slave_readdata                      (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),                   //                                                      .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                     (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),                  //                                                      .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                   (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest),                //                                                      .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                    (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),                 //                                                      .chipselect
		.nios2_gen2_0_debug_mem_slave_address                        (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address),                     //                          nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                          (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write),                       //                                                      .write
		.nios2_gen2_0_debug_mem_slave_read                           (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read),                        //                                                      .read
		.nios2_gen2_0_debug_mem_slave_readdata                       (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata),                    //                                                      .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                      (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata),                   //                                                      .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                     (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable),                  //                                                      .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                    (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest),                 //                                                      .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                    (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess),                 //                                                      .debugaccess
		.onchip_memory_s1_address                                    (mm_interconnect_1_onchip_memory_s1_address),                                 //                                      onchip_memory_s1.address
		.onchip_memory_s1_write                                      (mm_interconnect_1_onchip_memory_s1_write),                                   //                                                      .write
		.onchip_memory_s1_readdata                                   (mm_interconnect_1_onchip_memory_s1_readdata),                                //                                                      .readdata
		.onchip_memory_s1_writedata                                  (mm_interconnect_1_onchip_memory_s1_writedata),                               //                                                      .writedata
		.onchip_memory_s1_byteenable                                 (mm_interconnect_1_onchip_memory_s1_byteenable),                              //                                                      .byteenable
		.onchip_memory_s1_chipselect                                 (mm_interconnect_1_onchip_memory_s1_chipselect),                              //                                                      .chipselect
		.onchip_memory_s1_clken                                      (mm_interconnect_1_onchip_memory_s1_clken),                                   //                                                      .clken
		.rmap_mem_nfee_comm_1_avalon_rmap_slave_0_address            (mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_address),         //              rmap_mem_nfee_comm_1_avalon_rmap_slave_0.address
		.rmap_mem_nfee_comm_1_avalon_rmap_slave_0_write              (mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_write),           //                                                      .write
		.rmap_mem_nfee_comm_1_avalon_rmap_slave_0_read               (mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_read),            //                                                      .read
		.rmap_mem_nfee_comm_1_avalon_rmap_slave_0_readdata           (mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_readdata),        //                                                      .readdata
		.rmap_mem_nfee_comm_1_avalon_rmap_slave_0_writedata          (mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_writedata),       //                                                      .writedata
		.rmap_mem_nfee_comm_1_avalon_rmap_slave_0_byteenable         (mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_byteenable),      //                                                      .byteenable
		.rmap_mem_nfee_comm_1_avalon_rmap_slave_0_waitrequest        (mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_waitrequest),     //                                                      .waitrequest
		.rmap_mem_nfee_comm_2_avalon_rmap_slave_0_address            (mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_address),         //              rmap_mem_nfee_comm_2_avalon_rmap_slave_0.address
		.rmap_mem_nfee_comm_2_avalon_rmap_slave_0_write              (mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_write),           //                                                      .write
		.rmap_mem_nfee_comm_2_avalon_rmap_slave_0_read               (mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_read),            //                                                      .read
		.rmap_mem_nfee_comm_2_avalon_rmap_slave_0_readdata           (mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_readdata),        //                                                      .readdata
		.rmap_mem_nfee_comm_2_avalon_rmap_slave_0_writedata          (mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_writedata),       //                                                      .writedata
		.rmap_mem_nfee_comm_2_avalon_rmap_slave_0_byteenable         (mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_byteenable),      //                                                      .byteenable
		.rmap_mem_nfee_comm_2_avalon_rmap_slave_0_waitrequest        (mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_waitrequest),     //                                                      .waitrequest
		.rmap_mem_nfee_comm_3_avalon_rmap_slave_0_address            (mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_address),         //              rmap_mem_nfee_comm_3_avalon_rmap_slave_0.address
		.rmap_mem_nfee_comm_3_avalon_rmap_slave_0_write              (mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_write),           //                                                      .write
		.rmap_mem_nfee_comm_3_avalon_rmap_slave_0_read               (mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_read),            //                                                      .read
		.rmap_mem_nfee_comm_3_avalon_rmap_slave_0_readdata           (mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_readdata),        //                                                      .readdata
		.rmap_mem_nfee_comm_3_avalon_rmap_slave_0_writedata          (mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_writedata),       //                                                      .writedata
		.rmap_mem_nfee_comm_3_avalon_rmap_slave_0_byteenable         (mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_byteenable),      //                                                      .byteenable
		.rmap_mem_nfee_comm_3_avalon_rmap_slave_0_waitrequest        (mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_waitrequest),     //                                                      .waitrequest
		.rmap_mem_nfee_comm_4_avalon_rmap_slave_0_address            (mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_address),         //              rmap_mem_nfee_comm_4_avalon_rmap_slave_0.address
		.rmap_mem_nfee_comm_4_avalon_rmap_slave_0_write              (mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_write),           //                                                      .write
		.rmap_mem_nfee_comm_4_avalon_rmap_slave_0_read               (mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_read),            //                                                      .read
		.rmap_mem_nfee_comm_4_avalon_rmap_slave_0_readdata           (mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_readdata),        //                                                      .readdata
		.rmap_mem_nfee_comm_4_avalon_rmap_slave_0_writedata          (mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_writedata),       //                                                      .writedata
		.rmap_mem_nfee_comm_4_avalon_rmap_slave_0_byteenable         (mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_byteenable),      //                                                      .byteenable
		.rmap_mem_nfee_comm_4_avalon_rmap_slave_0_waitrequest        (mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_waitrequest),     //                                                      .waitrequest
		.rmap_mem_nfee_comm_5_avalon_rmap_slave_0_address            (mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_address),         //              rmap_mem_nfee_comm_5_avalon_rmap_slave_0.address
		.rmap_mem_nfee_comm_5_avalon_rmap_slave_0_write              (mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_write),           //                                                      .write
		.rmap_mem_nfee_comm_5_avalon_rmap_slave_0_read               (mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_read),            //                                                      .read
		.rmap_mem_nfee_comm_5_avalon_rmap_slave_0_readdata           (mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_readdata),        //                                                      .readdata
		.rmap_mem_nfee_comm_5_avalon_rmap_slave_0_writedata          (mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_writedata),       //                                                      .writedata
		.rmap_mem_nfee_comm_5_avalon_rmap_slave_0_byteenable         (mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_byteenable),      //                                                      .byteenable
		.rmap_mem_nfee_comm_5_avalon_rmap_slave_0_waitrequest        (mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_waitrequest),     //                                                      .waitrequest
		.rmap_mem_nfee_comm_6_avalon_rmap_slave_0_address            (mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_address),         //              rmap_mem_nfee_comm_6_avalon_rmap_slave_0.address
		.rmap_mem_nfee_comm_6_avalon_rmap_slave_0_write              (mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_write),           //                                                      .write
		.rmap_mem_nfee_comm_6_avalon_rmap_slave_0_read               (mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_read),            //                                                      .read
		.rmap_mem_nfee_comm_6_avalon_rmap_slave_0_readdata           (mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_readdata),        //                                                      .readdata
		.rmap_mem_nfee_comm_6_avalon_rmap_slave_0_writedata          (mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_writedata),       //                                                      .writedata
		.rmap_mem_nfee_comm_6_avalon_rmap_slave_0_byteenable         (mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_byteenable),      //                                                      .byteenable
		.rmap_mem_nfee_comm_6_avalon_rmap_slave_0_waitrequest        (mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_waitrequest),     //                                                      .waitrequest
		.sysid_qsys_control_slave_address                            (mm_interconnect_1_sysid_qsys_control_slave_address),                         //                              sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                           (mm_interconnect_1_sysid_qsys_control_slave_readdata)                         //                                                      .readdata
	);

	MebX_Qsys_Project_mm_interconnect_2 mm_interconnect_2 (
		.clk_50_clk_clk                                                         (clk50_clk),                                                                              //                                                       clk_50_clk.clk
		.Altera_UP_SD_Card_Avalon_Interface_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                                     // Altera_UP_SD_Card_Avalon_Interface_0_reset_reset_bridge_in_reset.reset
		.clock_bridge_afi_50_m0_reset_reset_bridge_in_reset_reset               (rst_controller_019_reset_out_reset),                                                     //               clock_bridge_afi_50_m0_reset_reset_bridge_in_reset.reset
		.rs232_uart_reset_reset_bridge_in_reset_reset                           (rst_controller_023_reset_out_reset),                                                     //                           rs232_uart_reset_reset_bridge_in_reset.reset
		.sync_reset_reset_bridge_in_reset_reset                                 (rst_controller_024_reset_out_reset),                                                     //                                 sync_reset_reset_bridge_in_reset.reset
		.clock_bridge_afi_50_m0_address                                         (clock_bridge_afi_50_m0_address),                                                         //                                           clock_bridge_afi_50_m0.address
		.clock_bridge_afi_50_m0_waitrequest                                     (clock_bridge_afi_50_m0_waitrequest),                                                     //                                                                 .waitrequest
		.clock_bridge_afi_50_m0_burstcount                                      (clock_bridge_afi_50_m0_burstcount),                                                      //                                                                 .burstcount
		.clock_bridge_afi_50_m0_byteenable                                      (clock_bridge_afi_50_m0_byteenable),                                                      //                                                                 .byteenable
		.clock_bridge_afi_50_m0_read                                            (clock_bridge_afi_50_m0_read),                                                            //                                                                 .read
		.clock_bridge_afi_50_m0_readdata                                        (clock_bridge_afi_50_m0_readdata),                                                        //                                                                 .readdata
		.clock_bridge_afi_50_m0_readdatavalid                                   (clock_bridge_afi_50_m0_readdatavalid),                                                   //                                                                 .readdatavalid
		.clock_bridge_afi_50_m0_write                                           (clock_bridge_afi_50_m0_write),                                                           //                                                                 .write
		.clock_bridge_afi_50_m0_writedata                                       (clock_bridge_afi_50_m0_writedata),                                                       //                                                                 .writedata
		.clock_bridge_afi_50_m0_debugaccess                                     (clock_bridge_afi_50_m0_debugaccess),                                                     //                                                                 .debugaccess
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address       (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address),     //         Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave.address
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write         (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write),       //                                                                 .write
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read          (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read),        //                                                                 .read
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata      (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata),    //                                                                 .readdata
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata     (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata),   //                                                                 .writedata
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable    (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable),  //                                                                 .byteenable
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest   (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest), //                                                                 .waitrequest
		.Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect    (mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect),  //                                                                 .chipselect
		.csense_adc_fo_s1_address                                               (mm_interconnect_2_csense_adc_fo_s1_address),                                             //                                                 csense_adc_fo_s1.address
		.csense_adc_fo_s1_write                                                 (mm_interconnect_2_csense_adc_fo_s1_write),                                               //                                                                 .write
		.csense_adc_fo_s1_readdata                                              (mm_interconnect_2_csense_adc_fo_s1_readdata),                                            //                                                                 .readdata
		.csense_adc_fo_s1_writedata                                             (mm_interconnect_2_csense_adc_fo_s1_writedata),                                           //                                                                 .writedata
		.csense_adc_fo_s1_chipselect                                            (mm_interconnect_2_csense_adc_fo_s1_chipselect),                                          //                                                                 .chipselect
		.csense_cs_n_s1_address                                                 (mm_interconnect_2_csense_cs_n_s1_address),                                               //                                                   csense_cs_n_s1.address
		.csense_cs_n_s1_write                                                   (mm_interconnect_2_csense_cs_n_s1_write),                                                 //                                                                 .write
		.csense_cs_n_s1_readdata                                                (mm_interconnect_2_csense_cs_n_s1_readdata),                                              //                                                                 .readdata
		.csense_cs_n_s1_writedata                                               (mm_interconnect_2_csense_cs_n_s1_writedata),                                             //                                                                 .writedata
		.csense_cs_n_s1_chipselect                                              (mm_interconnect_2_csense_cs_n_s1_chipselect),                                            //                                                                 .chipselect
		.csense_sck_s1_address                                                  (mm_interconnect_2_csense_sck_s1_address),                                                //                                                    csense_sck_s1.address
		.csense_sck_s1_write                                                    (mm_interconnect_2_csense_sck_s1_write),                                                  //                                                                 .write
		.csense_sck_s1_readdata                                                 (mm_interconnect_2_csense_sck_s1_readdata),                                               //                                                                 .readdata
		.csense_sck_s1_writedata                                                (mm_interconnect_2_csense_sck_s1_writedata),                                              //                                                                 .writedata
		.csense_sck_s1_chipselect                                               (mm_interconnect_2_csense_sck_s1_chipselect),                                             //                                                                 .chipselect
		.csense_sdi_s1_address                                                  (mm_interconnect_2_csense_sdi_s1_address),                                                //                                                    csense_sdi_s1.address
		.csense_sdi_s1_write                                                    (mm_interconnect_2_csense_sdi_s1_write),                                                  //                                                                 .write
		.csense_sdi_s1_readdata                                                 (mm_interconnect_2_csense_sdi_s1_readdata),                                               //                                                                 .readdata
		.csense_sdi_s1_writedata                                                (mm_interconnect_2_csense_sdi_s1_writedata),                                              //                                                                 .writedata
		.csense_sdi_s1_chipselect                                               (mm_interconnect_2_csense_sdi_s1_chipselect),                                             //                                                                 .chipselect
		.csense_sdo_s1_address                                                  (mm_interconnect_2_csense_sdo_s1_address),                                                //                                                    csense_sdo_s1.address
		.csense_sdo_s1_readdata                                                 (mm_interconnect_2_csense_sdo_s1_readdata),                                               //                                                                 .readdata
		.m1_ddr2_i2c_scl_s1_address                                             (mm_interconnect_2_m1_ddr2_i2c_scl_s1_address),                                           //                                               m1_ddr2_i2c_scl_s1.address
		.m1_ddr2_i2c_scl_s1_write                                               (mm_interconnect_2_m1_ddr2_i2c_scl_s1_write),                                             //                                                                 .write
		.m1_ddr2_i2c_scl_s1_readdata                                            (mm_interconnect_2_m1_ddr2_i2c_scl_s1_readdata),                                          //                                                                 .readdata
		.m1_ddr2_i2c_scl_s1_writedata                                           (mm_interconnect_2_m1_ddr2_i2c_scl_s1_writedata),                                         //                                                                 .writedata
		.m1_ddr2_i2c_scl_s1_chipselect                                          (mm_interconnect_2_m1_ddr2_i2c_scl_s1_chipselect),                                        //                                                                 .chipselect
		.m1_ddr2_i2c_sda_s1_address                                             (mm_interconnect_2_m1_ddr2_i2c_sda_s1_address),                                           //                                               m1_ddr2_i2c_sda_s1.address
		.m1_ddr2_i2c_sda_s1_write                                               (mm_interconnect_2_m1_ddr2_i2c_sda_s1_write),                                             //                                                                 .write
		.m1_ddr2_i2c_sda_s1_readdata                                            (mm_interconnect_2_m1_ddr2_i2c_sda_s1_readdata),                                          //                                                                 .readdata
		.m1_ddr2_i2c_sda_s1_writedata                                           (mm_interconnect_2_m1_ddr2_i2c_sda_s1_writedata),                                         //                                                                 .writedata
		.m1_ddr2_i2c_sda_s1_chipselect                                          (mm_interconnect_2_m1_ddr2_i2c_sda_s1_chipselect),                                        //                                                                 .chipselect
		.m2_ddr2_i2c_scl_s1_address                                             (mm_interconnect_2_m2_ddr2_i2c_scl_s1_address),                                           //                                               m2_ddr2_i2c_scl_s1.address
		.m2_ddr2_i2c_scl_s1_write                                               (mm_interconnect_2_m2_ddr2_i2c_scl_s1_write),                                             //                                                                 .write
		.m2_ddr2_i2c_scl_s1_readdata                                            (mm_interconnect_2_m2_ddr2_i2c_scl_s1_readdata),                                          //                                                                 .readdata
		.m2_ddr2_i2c_scl_s1_writedata                                           (mm_interconnect_2_m2_ddr2_i2c_scl_s1_writedata),                                         //                                                                 .writedata
		.m2_ddr2_i2c_scl_s1_chipselect                                          (mm_interconnect_2_m2_ddr2_i2c_scl_s1_chipselect),                                        //                                                                 .chipselect
		.m2_ddr2_i2c_sda_s1_address                                             (mm_interconnect_2_m2_ddr2_i2c_sda_s1_address),                                           //                                               m2_ddr2_i2c_sda_s1.address
		.m2_ddr2_i2c_sda_s1_write                                               (mm_interconnect_2_m2_ddr2_i2c_sda_s1_write),                                             //                                                                 .write
		.m2_ddr2_i2c_sda_s1_readdata                                            (mm_interconnect_2_m2_ddr2_i2c_sda_s1_readdata),                                          //                                                                 .readdata
		.m2_ddr2_i2c_sda_s1_writedata                                           (mm_interconnect_2_m2_ddr2_i2c_sda_s1_writedata),                                         //                                                                 .writedata
		.m2_ddr2_i2c_sda_s1_chipselect                                          (mm_interconnect_2_m2_ddr2_i2c_sda_s1_chipselect),                                        //                                                                 .chipselect
		.pio_BUTTON_s1_address                                                  (mm_interconnect_2_pio_button_s1_address),                                                //                                                    pio_BUTTON_s1.address
		.pio_BUTTON_s1_readdata                                                 (mm_interconnect_2_pio_button_s1_readdata),                                               //                                                                 .readdata
		.pio_ctrl_io_lvds_s1_address                                            (mm_interconnect_2_pio_ctrl_io_lvds_s1_address),                                          //                                              pio_ctrl_io_lvds_s1.address
		.pio_ctrl_io_lvds_s1_write                                              (mm_interconnect_2_pio_ctrl_io_lvds_s1_write),                                            //                                                                 .write
		.pio_ctrl_io_lvds_s1_readdata                                           (mm_interconnect_2_pio_ctrl_io_lvds_s1_readdata),                                         //                                                                 .readdata
		.pio_ctrl_io_lvds_s1_writedata                                          (mm_interconnect_2_pio_ctrl_io_lvds_s1_writedata),                                        //                                                                 .writedata
		.pio_ctrl_io_lvds_s1_chipselect                                         (mm_interconnect_2_pio_ctrl_io_lvds_s1_chipselect),                                       //                                                                 .chipselect
		.pio_DIP_s1_address                                                     (mm_interconnect_2_pio_dip_s1_address),                                                   //                                                       pio_DIP_s1.address
		.pio_DIP_s1_readdata                                                    (mm_interconnect_2_pio_dip_s1_readdata),                                                  //                                                                 .readdata
		.pio_EXT_s1_address                                                     (mm_interconnect_2_pio_ext_s1_address),                                                   //                                                       pio_EXT_s1.address
		.pio_EXT_s1_readdata                                                    (mm_interconnect_2_pio_ext_s1_readdata),                                                  //                                                                 .readdata
		.pio_LED_s1_address                                                     (mm_interconnect_2_pio_led_s1_address),                                                   //                                                       pio_LED_s1.address
		.pio_LED_s1_write                                                       (mm_interconnect_2_pio_led_s1_write),                                                     //                                                                 .write
		.pio_LED_s1_readdata                                                    (mm_interconnect_2_pio_led_s1_readdata),                                                  //                                                                 .readdata
		.pio_LED_s1_writedata                                                   (mm_interconnect_2_pio_led_s1_writedata),                                                 //                                                                 .writedata
		.pio_LED_s1_chipselect                                                  (mm_interconnect_2_pio_led_s1_chipselect),                                                //                                                                 .chipselect
		.pio_LED_painel_s1_address                                              (mm_interconnect_2_pio_led_painel_s1_address),                                            //                                                pio_LED_painel_s1.address
		.pio_LED_painel_s1_write                                                (mm_interconnect_2_pio_led_painel_s1_write),                                              //                                                                 .write
		.pio_LED_painel_s1_readdata                                             (mm_interconnect_2_pio_led_painel_s1_readdata),                                           //                                                                 .readdata
		.pio_LED_painel_s1_writedata                                            (mm_interconnect_2_pio_led_painel_s1_writedata),                                          //                                                                 .writedata
		.pio_LED_painel_s1_chipselect                                           (mm_interconnect_2_pio_led_painel_s1_chipselect),                                         //                                                                 .chipselect
		.rs232_uart_s1_address                                                  (mm_interconnect_2_rs232_uart_s1_address),                                                //                                                    rs232_uart_s1.address
		.rs232_uart_s1_write                                                    (mm_interconnect_2_rs232_uart_s1_write),                                                  //                                                                 .write
		.rs232_uart_s1_read                                                     (mm_interconnect_2_rs232_uart_s1_read),                                                   //                                                                 .read
		.rs232_uart_s1_readdata                                                 (mm_interconnect_2_rs232_uart_s1_readdata),                                               //                                                                 .readdata
		.rs232_uart_s1_writedata                                                (mm_interconnect_2_rs232_uart_s1_writedata),                                              //                                                                 .writedata
		.rs232_uart_s1_begintransfer                                            (mm_interconnect_2_rs232_uart_s1_begintransfer),                                          //                                                                 .begintransfer
		.rs232_uart_s1_chipselect                                               (mm_interconnect_2_rs232_uart_s1_chipselect),                                             //                                                                 .chipselect
		.rst_controller_avalon_rst_controller_slave_address                     (mm_interconnect_2_rst_controller_avalon_rst_controller_slave_address),                   //                       rst_controller_avalon_rst_controller_slave.address
		.rst_controller_avalon_rst_controller_slave_write                       (mm_interconnect_2_rst_controller_avalon_rst_controller_slave_write),                     //                                                                 .write
		.rst_controller_avalon_rst_controller_slave_read                        (mm_interconnect_2_rst_controller_avalon_rst_controller_slave_read),                      //                                                                 .read
		.rst_controller_avalon_rst_controller_slave_readdata                    (mm_interconnect_2_rst_controller_avalon_rst_controller_slave_readdata),                  //                                                                 .readdata
		.rst_controller_avalon_rst_controller_slave_writedata                   (mm_interconnect_2_rst_controller_avalon_rst_controller_slave_writedata),                 //                                                                 .writedata
		.rst_controller_avalon_rst_controller_slave_waitrequest                 (mm_interconnect_2_rst_controller_avalon_rst_controller_slave_waitrequest),               //                                                                 .waitrequest
		.rtcc_alarm_s1_address                                                  (mm_interconnect_2_rtcc_alarm_s1_address),                                                //                                                    rtcc_alarm_s1.address
		.rtcc_alarm_s1_readdata                                                 (mm_interconnect_2_rtcc_alarm_s1_readdata),                                               //                                                                 .readdata
		.rtcc_cs_n_s1_address                                                   (mm_interconnect_2_rtcc_cs_n_s1_address),                                                 //                                                     rtcc_cs_n_s1.address
		.rtcc_cs_n_s1_write                                                     (mm_interconnect_2_rtcc_cs_n_s1_write),                                                   //                                                                 .write
		.rtcc_cs_n_s1_readdata                                                  (mm_interconnect_2_rtcc_cs_n_s1_readdata),                                                //                                                                 .readdata
		.rtcc_cs_n_s1_writedata                                                 (mm_interconnect_2_rtcc_cs_n_s1_writedata),                                               //                                                                 .writedata
		.rtcc_cs_n_s1_chipselect                                                (mm_interconnect_2_rtcc_cs_n_s1_chipselect),                                              //                                                                 .chipselect
		.rtcc_sck_s1_address                                                    (mm_interconnect_2_rtcc_sck_s1_address),                                                  //                                                      rtcc_sck_s1.address
		.rtcc_sck_s1_write                                                      (mm_interconnect_2_rtcc_sck_s1_write),                                                    //                                                                 .write
		.rtcc_sck_s1_readdata                                                   (mm_interconnect_2_rtcc_sck_s1_readdata),                                                 //                                                                 .readdata
		.rtcc_sck_s1_writedata                                                  (mm_interconnect_2_rtcc_sck_s1_writedata),                                                //                                                                 .writedata
		.rtcc_sck_s1_chipselect                                                 (mm_interconnect_2_rtcc_sck_s1_chipselect),                                               //                                                                 .chipselect
		.rtcc_sdi_s1_address                                                    (mm_interconnect_2_rtcc_sdi_s1_address),                                                  //                                                      rtcc_sdi_s1.address
		.rtcc_sdi_s1_write                                                      (mm_interconnect_2_rtcc_sdi_s1_write),                                                    //                                                                 .write
		.rtcc_sdi_s1_readdata                                                   (mm_interconnect_2_rtcc_sdi_s1_readdata),                                                 //                                                                 .readdata
		.rtcc_sdi_s1_writedata                                                  (mm_interconnect_2_rtcc_sdi_s1_writedata),                                                //                                                                 .writedata
		.rtcc_sdi_s1_chipselect                                                 (mm_interconnect_2_rtcc_sdi_s1_chipselect),                                               //                                                                 .chipselect
		.rtcc_sdo_s1_address                                                    (mm_interconnect_2_rtcc_sdo_s1_address),                                                  //                                                      rtcc_sdo_s1.address
		.rtcc_sdo_s1_readdata                                                   (mm_interconnect_2_rtcc_sdo_s1_readdata),                                                 //                                                                 .readdata
		.sd_card_wp_n_s1_address                                                (mm_interconnect_2_sd_card_wp_n_s1_address),                                              //                                                  sd_card_wp_n_s1.address
		.sd_card_wp_n_s1_readdata                                               (mm_interconnect_2_sd_card_wp_n_s1_readdata),                                             //                                                                 .readdata
		.sync_avalon_mm_slave_address                                           (mm_interconnect_2_sync_avalon_mm_slave_address),                                         //                                             sync_avalon_mm_slave.address
		.sync_avalon_mm_slave_write                                             (mm_interconnect_2_sync_avalon_mm_slave_write),                                           //                                                                 .write
		.sync_avalon_mm_slave_read                                              (mm_interconnect_2_sync_avalon_mm_slave_read),                                            //                                                                 .read
		.sync_avalon_mm_slave_readdata                                          (mm_interconnect_2_sync_avalon_mm_slave_readdata),                                        //                                                                 .readdata
		.sync_avalon_mm_slave_writedata                                         (mm_interconnect_2_sync_avalon_mm_slave_writedata),                                       //                                                                 .writedata
		.sync_avalon_mm_slave_byteenable                                        (mm_interconnect_2_sync_avalon_mm_slave_byteenable),                                      //                                                                 .byteenable
		.sync_avalon_mm_slave_waitrequest                                       (mm_interconnect_2_sync_avalon_mm_slave_waitrequest),                                     //                                                                 .waitrequest
		.temp_scl_s1_address                                                    (mm_interconnect_2_temp_scl_s1_address),                                                  //                                                      temp_scl_s1.address
		.temp_scl_s1_write                                                      (mm_interconnect_2_temp_scl_s1_write),                                                    //                                                                 .write
		.temp_scl_s1_readdata                                                   (mm_interconnect_2_temp_scl_s1_readdata),                                                 //                                                                 .readdata
		.temp_scl_s1_writedata                                                  (mm_interconnect_2_temp_scl_s1_writedata),                                                //                                                                 .writedata
		.temp_scl_s1_chipselect                                                 (mm_interconnect_2_temp_scl_s1_chipselect),                                               //                                                                 .chipselect
		.temp_sda_s1_address                                                    (mm_interconnect_2_temp_sda_s1_address),                                                  //                                                      temp_sda_s1.address
		.temp_sda_s1_write                                                      (mm_interconnect_2_temp_sda_s1_write),                                                    //                                                                 .write
		.temp_sda_s1_readdata                                                   (mm_interconnect_2_temp_sda_s1_readdata),                                                 //                                                                 .readdata
		.temp_sda_s1_writedata                                                  (mm_interconnect_2_temp_sda_s1_writedata),                                                //                                                                 .writedata
		.temp_sda_s1_chipselect                                                 (mm_interconnect_2_temp_sda_s1_chipselect),                                               //                                                                 .chipselect
		.timer_1ms_s1_address                                                   (mm_interconnect_2_timer_1ms_s1_address),                                                 //                                                     timer_1ms_s1.address
		.timer_1ms_s1_write                                                     (mm_interconnect_2_timer_1ms_s1_write),                                                   //                                                                 .write
		.timer_1ms_s1_readdata                                                  (mm_interconnect_2_timer_1ms_s1_readdata),                                                //                                                                 .readdata
		.timer_1ms_s1_writedata                                                 (mm_interconnect_2_timer_1ms_s1_writedata),                                               //                                                                 .writedata
		.timer_1ms_s1_chipselect                                                (mm_interconnect_2_timer_1ms_s1_chipselect),                                              //                                                                 .chipselect
		.timer_1us_s1_address                                                   (mm_interconnect_2_timer_1us_s1_address),                                                 //                                                     timer_1us_s1.address
		.timer_1us_s1_write                                                     (mm_interconnect_2_timer_1us_s1_write),                                                   //                                                                 .write
		.timer_1us_s1_readdata                                                  (mm_interconnect_2_timer_1us_s1_readdata),                                                //                                                                 .readdata
		.timer_1us_s1_writedata                                                 (mm_interconnect_2_timer_1us_s1_writedata),                                               //                                                                 .writedata
		.timer_1us_s1_chipselect                                                (mm_interconnect_2_timer_1us_s1_chipselect)                                               //                                                                 .chipselect
	);

	MebX_Qsys_Project_mm_interconnect_3 mm_interconnect_3 (
		.m1_ddr2_memory_afi_clk_clk                                      (m1_ddr2_memory_afi_clk_clk),                              //                                    m1_ddr2_memory_afi_clk.clk
		.m1_ddr2_memory_afi_half_clk_clk                                 (m1_ddr2_memory_afi_half_clk_clk),                         //                               m1_ddr2_memory_afi_half_clk.clk
		.m1_clock_bridge_m0_reset_reset_bridge_in_reset_reset            (rst_controller_021_reset_out_reset),                      //            m1_clock_bridge_m0_reset_reset_bridge_in_reset.reset
		.m1_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset (rst_controller_026_reset_out_reset),                      // m1_ddr2_memory_avl_translator_reset_reset_bridge_in_reset.reset
		.m1_ddr2_memory_soft_reset_reset_bridge_in_reset_reset           (rst_controller_026_reset_out_reset),                      //           m1_ddr2_memory_soft_reset_reset_bridge_in_reset.reset
		.m1_clock_bridge_m0_address                                      (m1_clock_bridge_m0_address),                              //                                        m1_clock_bridge_m0.address
		.m1_clock_bridge_m0_waitrequest                                  (m1_clock_bridge_m0_waitrequest),                          //                                                          .waitrequest
		.m1_clock_bridge_m0_burstcount                                   (m1_clock_bridge_m0_burstcount),                           //                                                          .burstcount
		.m1_clock_bridge_m0_byteenable                                   (m1_clock_bridge_m0_byteenable),                           //                                                          .byteenable
		.m1_clock_bridge_m0_read                                         (m1_clock_bridge_m0_read),                                 //                                                          .read
		.m1_clock_bridge_m0_readdata                                     (m1_clock_bridge_m0_readdata),                             //                                                          .readdata
		.m1_clock_bridge_m0_readdatavalid                                (m1_clock_bridge_m0_readdatavalid),                        //                                                          .readdatavalid
		.m1_clock_bridge_m0_write                                        (m1_clock_bridge_m0_write),                                //                                                          .write
		.m1_clock_bridge_m0_writedata                                    (m1_clock_bridge_m0_writedata),                            //                                                          .writedata
		.m1_clock_bridge_m0_debugaccess                                  (m1_clock_bridge_m0_debugaccess),                          //                                                          .debugaccess
		.m1_ddr2_memory_avl_address                                      (mm_interconnect_3_m1_ddr2_memory_avl_address),            //                                        m1_ddr2_memory_avl.address
		.m1_ddr2_memory_avl_write                                        (mm_interconnect_3_m1_ddr2_memory_avl_write),              //                                                          .write
		.m1_ddr2_memory_avl_read                                         (mm_interconnect_3_m1_ddr2_memory_avl_read),               //                                                          .read
		.m1_ddr2_memory_avl_readdata                                     (mm_interconnect_3_m1_ddr2_memory_avl_readdata),           //                                                          .readdata
		.m1_ddr2_memory_avl_writedata                                    (mm_interconnect_3_m1_ddr2_memory_avl_writedata),          //                                                          .writedata
		.m1_ddr2_memory_avl_beginbursttransfer                           (mm_interconnect_3_m1_ddr2_memory_avl_beginbursttransfer), //                                                          .beginbursttransfer
		.m1_ddr2_memory_avl_burstcount                                   (mm_interconnect_3_m1_ddr2_memory_avl_burstcount),         //                                                          .burstcount
		.m1_ddr2_memory_avl_byteenable                                   (mm_interconnect_3_m1_ddr2_memory_avl_byteenable),         //                                                          .byteenable
		.m1_ddr2_memory_avl_readdatavalid                                (mm_interconnect_3_m1_ddr2_memory_avl_readdatavalid),      //                                                          .readdatavalid
		.m1_ddr2_memory_avl_waitrequest                                  (~mm_interconnect_3_m1_ddr2_memory_avl_waitrequest)        //                                                          .waitrequest
	);

	MebX_Qsys_Project_irq_mapper irq_mapper (
		.clk            (m2_ddr2_memory_afi_half_clk_clk),    //        clk.clk
		.reset          (rst_controller_022_reset_out_reset), //  clk_reset.reset
		.receiver0_irq  (irq_mapper_receiver0_irq),           //  receiver0.irq
		.receiver1_irq  (irq_mapper_receiver1_irq),           //  receiver1.irq
		.receiver2_irq  (irq_mapper_receiver2_irq),           //  receiver2.irq
		.receiver3_irq  (irq_mapper_receiver3_irq),           //  receiver3.irq
		.receiver4_irq  (irq_mapper_receiver4_irq),           //  receiver4.irq
		.receiver5_irq  (irq_mapper_receiver5_irq),           //  receiver5.irq
		.receiver6_irq  (irq_mapper_receiver6_irq),           //  receiver6.irq
		.receiver7_irq  (irq_mapper_receiver7_irq),           //  receiver7.irq
		.receiver8_irq  (irq_mapper_receiver8_irq),           //  receiver8.irq
		.receiver9_irq  (irq_mapper_receiver9_irq),           //  receiver9.irq
		.receiver10_irq (irq_mapper_receiver10_irq),          // receiver10.irq
		.receiver11_irq (irq_mapper_receiver11_irq),          // receiver11.irq
		.receiver12_irq (irq_mapper_receiver12_irq),          // receiver12.irq
		.receiver13_irq (irq_mapper_receiver13_irq),          // receiver13.irq
		.receiver14_irq (irq_mapper_receiver14_irq),          // receiver14.irq
		.receiver15_irq (irq_mapper_receiver15_irq),          // receiver15.irq
		.receiver16_irq (irq_mapper_receiver16_irq),          // receiver16.irq
		.receiver17_irq (irq_mapper_receiver17_irq),          // receiver17.irq
		.receiver18_irq (irq_mapper_receiver18_irq),          // receiver18.irq
		.receiver19_irq (irq_mapper_receiver19_irq),          // receiver19.irq
		.sender_irq     (nios2_gen2_0_irq_irq)                //     sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk50_clk),                          //       receiver_clk.clk
		.sender_clk     (m2_ddr2_memory_afi_half_clk_clk),    //         sender_clk.clk
		.receiver_reset (rst_controller_019_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_022_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver9_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk50_clk),                          //       receiver_clk.clk
		.sender_clk     (m2_ddr2_memory_afi_half_clk_clk),    //         sender_clk.clk
		.receiver_reset (rst_controller_019_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_022_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver10_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk50_clk),                          //       receiver_clk.clk
		.sender_clk     (m2_ddr2_memory_afi_half_clk_clk),    //         sender_clk.clk
		.receiver_reset (rst_controller_023_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_022_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver11_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk50_clk),                          //       receiver_clk.clk
		.sender_clk     (m2_ddr2_memory_afi_half_clk_clk),    //         sender_clk.clk
		.receiver_reset (rst_controller_024_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_022_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver12_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (clk50_clk),                          //       receiver_clk.clk
		.sender_clk     (m2_ddr2_memory_afi_half_clk_clk),    //         sender_clk.clk
		.receiver_reset (rst_controller_024_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_022_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver19_irq)           //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~rst_reset_n),                              // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_sd_card_reset), // reset_in1.reset
		.clk            (clk50_clk),                                 //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),        // reset_out.reset
		.reset_req      (),                                          // (terminated)
		.reset_req_in0  (1'b0),                                      // (terminated)
		.reset_req_in1  (1'b0),                                      // (terminated)
		.reset_in2      (1'b0),                                      // (terminated)
		.reset_req_in2  (1'b0),                                      // (terminated)
		.reset_in3      (1'b0),                                      // (terminated)
		.reset_req_in3  (1'b0),                                      // (terminated)
		.reset_in4      (1'b0),                                      // (terminated)
		.reset_req_in4  (1'b0),                                      // (terminated)
		.reset_in5      (1'b0),                                      // (terminated)
		.reset_req_in5  (1'b0),                                      // (terminated)
		.reset_in6      (1'b0),                                      // (terminated)
		.reset_req_in6  (1'b0),                                      // (terminated)
		.reset_in7      (1'b0),                                      // (terminated)
		.reset_req_in7  (1'b0),                                      // (terminated)
		.reset_in8      (1'b0),                                      // (terminated)
		.reset_req_in8  (1'b0),                                      // (terminated)
		.reset_in9      (1'b0),                                      // (terminated)
		.reset_req_in9  (1'b0),                                      // (terminated)
		.reset_in10     (1'b0),                                      // (terminated)
		.reset_req_in10 (1'b0),                                      // (terminated)
		.reset_in11     (1'b0),                                      // (terminated)
		.reset_req_in11 (1'b0),                                      // (terminated)
		.reset_in12     (1'b0),                                      // (terminated)
		.reset_req_in12 (1'b0),                                      // (terminated)
		.reset_in13     (1'b0),                                      // (terminated)
		.reset_req_in13 (1'b0),                                      // (terminated)
		.reset_in14     (1'b0),                                      // (terminated)
		.reset_req_in14 (1'b0),                                      // (terminated)
		.reset_in15     (1'b0),                                      // (terminated)
		.reset_req_in15 (1'b0)                                       // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch1_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_half_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch2_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_half_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch3_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_half_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch4_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_half_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch5_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_half_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_007 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch6_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_half_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_007_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_008 (
		.reset_in0      (~rst_reset_n),                           // reset_in0.reset
		.clk            (m2_ddr2_memory_afi_half_clk_clk),        //       clk.clk
		.reset_out      (rst_controller_008_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_008_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (9),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_009 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch1_reset), // reset_in1.reset
		.reset_in2      (rst_controller_reset_source_comm_ch2_reset), // reset_in2.reset
		.reset_in3      (rst_controller_reset_source_comm_ch3_reset), // reset_in3.reset
		.reset_in4      (rst_controller_reset_source_comm_ch4_reset), // reset_in4.reset
		.reset_in5      (rst_controller_reset_source_comm_ch5_reset), // reset_in5.reset
		.reset_in6      (rst_controller_reset_source_comm_ch6_reset), // reset_in6.reset
		.reset_in7      (rst_controller_reset_source_comm_ch7_reset), // reset_in7.reset
		.reset_in8      (rst_controller_reset_source_comm_ch8_reset), // reset_in8.reset
		.clk            (m2_ddr2_memory_afi_half_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_009_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_010 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch1_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_010_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_011 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch2_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_011_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_012 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch3_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_012_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_013 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch4_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_013_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_014 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch5_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_014_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_015 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch6_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_015_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_016 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch7_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_016_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_017 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch8_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_017_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_018 (
		.reset_in0      (~rst_reset_n),                               // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_comm_ch7_reset), // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_half_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_018_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_019 (
		.reset_in0      (~rst_reset_n),                       // reset_in0.reset
		.clk            (clk50_clk),                          //       clk.clk
		.reset_out      (rst_controller_019_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_020 (
		.reset_in0      (~rst_reset_n),                       // reset_in0.reset
		.reset_in1      (~rst_reset_n),                       // reset_in1.reset
		.clk            (m2_ddr2_memory_afi_half_clk_clk),    //       clk.clk
		.reset_out      (rst_controller_020_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_021 (
		.reset_in0      (~rst_reset_n),                       // reset_in0.reset
		.clk            (m1_ddr2_memory_afi_half_clk_clk),    //       clk.clk
		.reset_out      (rst_controller_021_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_022 (
		.reset_in0      (~rst_reset_n),                           // reset_in0.reset
		.clk            (m2_ddr2_memory_afi_half_clk_clk),        //       clk.clk
		.reset_out      (rst_controller_022_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_022_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_023 (
		.reset_in0      (~rst_reset_n),                            // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_rs232_reset), // reset_in1.reset
		.clk            (clk50_clk),                               //       clk.clk
		.reset_out      (rst_controller_023_reset_out_reset),      // reset_out.reset
		.reset_req      (),                                        // (terminated)
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_024 (
		.reset_in0      (~rst_reset_n),                           // reset_in0.reset
		.reset_in1      (rst_controller_reset_source_sync_reset), // reset_in1.reset
		.clk            (clk50_clk),                              //       clk.clk
		.reset_out      (rst_controller_024_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_025 (
		.reset_in0      (~rst_reset_n),                       // reset_in0.reset
		.clk            (m2_ddr2_memory_afi_clk_clk),         //       clk.clk
		.reset_out      (rst_controller_025_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_026 (
		.reset_in0      (~rst_reset_n),                       // reset_in0.reset
		.clk            (m1_ddr2_memory_afi_clk_clk),         //       clk.clk
		.reset_out      (rst_controller_026_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
