package rmap_target_registers_pkg is
	
end package rmap_target_registers_pkg;

package body rmap_target_registers_pkg is
	
end package body rmap_target_registers_pkg;
