package rmap_target_write_reply_header_header_crc_pkg is
	
end package rmap_target_write_reply_header_header_crc_pkg;

package body rmap_target_write_reply_header_header_crc_pkg is
	
end package body rmap_target_write_reply_header_header_crc_pkg;
