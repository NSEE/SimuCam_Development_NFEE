--N�cleo de Sistemas Embarcados - Instituto Mau� de Tecnologia
--projeto: Simulador FEE
--nome do programa: 
--finalidade: Finalidade do programa
--vers�o: 1.0
--autor: Tiago Sanches da Silva
--                 <tiago.eem@gmail.com>
--data: 01-09-11
-------------------------------------------------------------------------------
--Modify : 25/09 - Rafael Corsi
--
-- Data and control to falling edge
-------------------------------------------------------------------------------
-- ======================
-- Modificacoes - Corsi
-- ======================
-- PLATO 2.0 - set/2014
-------------------------------------------------------------------------------
-- removido atualizacao do valor em borda de decida, isso implica em melhor
-- desempenho. 
-- Removido registradores extras colocado quando os sianis eram alterados em 
-- borda de subida
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity GlobalMux is
  port
    (

      clock                : in std_logic;
      Sel_DMux_nWrite_Data : in std_logic_vector(2 downto 0);  -- (000:Head;001:DataBody;010:HK;011:Read; 1XX: EEP)

      nWrite_Head     : in std_logic;
      nWrite_DataBody : in std_logic;
      nWrite_Read     : in std_logic;
      nWrite_Control  : in std_logic;

      data_Head     : in std_logic_vector(8 downto 0);
      data_DataBody : in std_logic_vector(8 downto 0);
      data_Read     : in std_logic_vector(8 downto 0);

      nWrite_out : out std_logic;
      data_out   : out std_logic_vector(8 downto 0)

      );

end GlobalMux;

architecture rtl of GlobalMux is

  signal nWrite_int : std_logic := '1';
  signal data_int   : std_logic_vector(8 downto 0) := (others => '0') ;
    
begin

  process(Sel_DMux_nWrite_Data, data_Head, nWrite_Head, 
			data_DataBody, nWrite_DataBody, 	
			data_Read, nWrite_Read,
			nWrite_Control)
  begin
      case Sel_DMux_nWrite_Data is
        when "000" =>
          data_int   <= data_Head;
          nWrite_int <= nWrite_Head;
        when "001" =>
          data_int   <= data_DataBody;
          nWrite_int <= nWrite_DataBody;
        when "011" =>
          data_int   <= data_Read;
          nWrite_int <= nWrite_Read;
        when others =>                  --eep
          data_int <= "100000001";
          nWrite_int <= nWrite_Control; -- error generated by controller
      end case;
  end process;

  data_out   <= data_int;
  nwrite_out <= nWrite_int;

    
end rtl;





