library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fee_data_controller_top is
	port(
		clk_i : in std_logic;
		rst_i : in std_logic
	);
end entity fee_data_controller_top;

architecture RTL of fee_data_controller_top is

begin

end architecture RTL;
