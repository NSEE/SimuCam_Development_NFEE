TX_LVDS_inst : TX_LVDS PORT MAP (
		tx_in	 => tx_in_sig,
		tx_out	 => tx_out_sig
	);
