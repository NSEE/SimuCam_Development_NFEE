library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity avalon_stimuli is
	port(
		clk : in std_logic;
		rst : in std_logic
	);
end entity avalon_stimuli;

architecture RTL of avalon_stimuli is
	
begin

end architecture RTL;
