package rmap_target_read_pkg is
	
end package rmap_target_read_pkg;

package body rmap_target_read_pkg is
	
end package body rmap_target_read_pkg;
