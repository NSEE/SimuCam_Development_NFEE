spwr_dvriso_en_out_altiobuf_inst : spwr_dvriso_en_out_altiobuf PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig
	);
