package rmap_target_pkg is
	
end package rmap_target_pkg;

package body rmap_target_pkg is
	
end package body rmap_target_pkg;
