package rmap_target_read_reply_header_data_length_pkg is
	
end package rmap_target_read_reply_header_data_length_pkg;

package body rmap_target_read_reply_header_data_length_pkg is
	
end package body rmap_target_read_reply_header_data_length_pkg;
