library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ftdi_data_receiver_ent is
	port(
		clk_i : in std_logic;
		rst_i : in std_logic
	);
end entity ftdi_data_receiver_ent;

architecture RTL of ftdi_data_receiver_ent is
	
begin

end architecture RTL;
