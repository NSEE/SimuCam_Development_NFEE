library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sync_outmux_ent is
	port(
		clk_i : in std_logic;
		rst_i : in std_logic
	);
end entity sync_outmux_ent;

architecture RTL of sync_outmux_ent is
	
begin

end architecture RTL;
