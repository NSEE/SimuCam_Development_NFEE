package rmap_target_write_reply_header_eop_pkg is
	
end package rmap_target_write_reply_header_eop_pkg;

package body rmap_target_write_reply_header_eop_pkg is
	
end package body rmap_target_write_reply_header_eop_pkg;
