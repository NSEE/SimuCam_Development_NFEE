-- megafunction wizard: %ALTIOBUF%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altiobuf_in 

-- ============================================================
-- File Name: spwr_select_in_altiobuf.vhd
-- Megafunction Name(s):
-- 			altiobuf_in
--
-- Simulation Library Files(s):
-- 			stratixiv
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Standard Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


--altiobuf_in CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" ENABLE_BUS_HOLD="FALSE" NUMBER_OF_CHANNELS=2 USE_DIFFERENTIAL_MODE="FALSE" USE_DYNAMIC_TERMINATION_CONTROL="FALSE" datain dataout
--VERSION_BEGIN 18.1 cbx_altiobuf_in 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_stratixiii 2018:09:12:13:04:24:SJ cbx_stratixv 2018:09:12:13:04:24:SJ  VERSION_END

 LIBRARY stratixiv;
 USE stratixiv.all;

--synthesis_resources = stratixiv_io_ibuf 2 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  spwr_select_in_altiobuf_iobuf_in_b5i IS 
	 PORT 
	 ( 
		 datain	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 dataout	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	 ); 
 END spwr_select_in_altiobuf_iobuf_in_b5i;

 ARCHITECTURE RTL OF spwr_select_in_altiobuf_iobuf_in_b5i IS

	 SIGNAL  wire_ibufa_i	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_ibufa_o	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 COMPONENT  stratixiv_io_ibuf
	 GENERIC 
	 (
		bus_hold	:	STRING := "false";
		differential_mode	:	STRING := "false";
		simulate_z_as	:	STRING := "Z";
		lpm_type	:	STRING := "stratixiv_io_ibuf"
	 );
	 PORT
	 ( 
		dynamicterminationcontrol	:	IN STD_LOGIC := '0';
		i	:	IN STD_LOGIC := '0';
		ibar	:	IN STD_LOGIC := '0';
		o	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	dataout <= wire_ibufa_o;
	wire_ibufa_i <= datain;
	loop0 : FOR i IN 0 TO 1 GENERATE 
	  ibufa :  stratixiv_io_ibuf
	  GENERIC MAP (
		bus_hold => "false",
		differential_mode => "false"
	  )
	  PORT MAP ( 
		i => wire_ibufa_i(i),
		o => wire_ibufa_o(i)
	  );
	END GENERATE loop0;

 END RTL; --spwr_select_in_altiobuf_iobuf_in_b5i
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY spwr_select_in_altiobuf IS
	PORT
	(
		datain		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		dataout		: OUT STD_LOGIC_VECTOR (1 DOWNTO 0)
	);
END spwr_select_in_altiobuf;


ARCHITECTURE RTL OF spwr_select_in_altiobuf IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (1 DOWNTO 0);



	COMPONENT spwr_select_in_altiobuf_iobuf_in_b5i
	PORT (
			datain	: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
			dataout	: OUT STD_LOGIC_VECTOR (1 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	dataout    <= sub_wire0(1 DOWNTO 0);

	spwr_select_in_altiobuf_iobuf_in_b5i_component : spwr_select_in_altiobuf_iobuf_in_b5i
	PORT MAP (
		datain => datain,
		dataout => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "1"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
-- Retrieval info: CONSTANT: enable_bus_hold STRING "FALSE"
-- Retrieval info: CONSTANT: number_of_channels NUMERIC "2"
-- Retrieval info: CONSTANT: use_differential_mode STRING "FALSE"
-- Retrieval info: CONSTANT: use_dynamic_termination_control STRING "FALSE"
-- Retrieval info: USED_PORT: datain 0 0 2 0 INPUT NODEFVAL "datain[1..0]"
-- Retrieval info: USED_PORT: dataout 0 0 2 0 OUTPUT NODEFVAL "dataout[1..0]"
-- Retrieval info: CONNECT: @datain 0 0 2 0 datain 0 0 2 0
-- Retrieval info: CONNECT: dataout 0 0 2 0 @dataout 0 0 2 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL spwr_select_in_altiobuf.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL spwr_select_in_altiobuf.inc TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL spwr_select_in_altiobuf.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL spwr_select_in_altiobuf.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL spwr_select_in_altiobuf_inst.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL spwr_select_in_altiobuf_syn.v TRUE
-- Retrieval info: LIB_FILE: stratixiv
