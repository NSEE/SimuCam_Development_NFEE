spwc_leds_out_altiobuf_inst : spwc_leds_out_altiobuf PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig
	);
