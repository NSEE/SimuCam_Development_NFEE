io_inout_39b_inst : io_inout_39b PORT MAP (
		datain	 => datain_sig,
		oe	 => oe_sig,
		dataio	 => dataio_sig,
		dataout	 => dataout_sig
	);
