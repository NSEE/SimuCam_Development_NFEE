package package is
	
end package package;

package body package is
	
end package body package;
