spwc_spw_tx_altiobuf_inst : spwc_spw_tx_altiobuf PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig,
		dataout_b	 => dataout_b_sig
	);
