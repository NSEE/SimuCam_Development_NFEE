// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
APztJhjEx1DJiMgJYytwbnQE46vd6APYAJ8VuAfwXELsei3jj+dC8U4UJz3g7PPpZyyOV5DREOZo
ouomBAE0DaYB0xQARC6mpDurqnX1uDmlL0ac+MGnv36FiUb1z1w7yLGDOgjoSap5h2Sv33SFHTfP
2PyFQZaT7BJlTy2zYqppQBcOaSrQ4nRUSvI2q9Qf2j8CZ9f4NCrl+q+2nn41GXCZETFKGcpizDbL
h2Y5ospP1ZdUAYqucpcOCgczNqV1cjZ7eg5APWSJM1Ws20q+1OwnO7T1Z47AxdFHh3E3Axl8vXAf
0/sZ1eXmCGHiwZfYONH+EEhp8QcNaNszkxFQcw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 16912)
OFwmtXArWC/wTQ+3sImwFCMf9Pj1RomFKJClK8O67uazE21+oFWd07WnRP48pa0eAruHQ85W7b0f
RHQF8aY84rQSKessd/7gIBqwnkdHpQ60Z87ncT0RtAQzllU5ouxrngz4mlrbFAQGYkHBGdfn5oDf
M9sNxgshwcz028jL/8eKNcjO/JJ1xJ2HMBNQ6ooAedAxHaoF2YJaGfPNU2xM8pmDbuhPvk//stvg
qwQnEf5bYOISJWsvLbJB6FnMFUlakROzjztw0F24Dpsd/bPTZfMvrBBJyGoLkdEYOaQXiyepocf5
e96MPHVg7xQVnIc3nEPdHeRUyxXNRC4mVAKI2aO0Oxpw3HQwIYjb/dm6U+Zv/GK7NkiQdXxgupox
+4LCmZaOEoHCHHmJgIb8JLHRfnTg8s9t31s4nOx2xloOeadfqXzmh5SBTJBtWomKPKNYH2VDeyJY
qeoQtq2JRHr0XwO2AMcb3eZ5GLgDKdUYpva4NICZaM18XNjAyCthjIujtPamU57jgZVNomHlG43m
m1ggO3Mp1gvHzfGtWYQFZwcpeLCzeSlAtDt5RWJNF0sdLI9/bkGwHaZrEKyFZjAdw9atk4toAU+T
ZcdUnFoxTTSYbprt/xbNAneiMB2YQRJxPGhhNLDDDTanB2LZQZrmuGMxB1c0XATuioXCzVG9gW7v
sJut0jUQiWgCf6+2YuAbe+M81T8hku0PeqmaG8N4E1Y4doPQFRRhXxLFns/zHF619Z+l9s+Ta4w6
MyAhqkZbLF7XRwSbgBeRzYi0nJEmSG2D+hKAmJP1xN7+6mvrtPeNgNyt715N5RrSbMJv0rfDX8Ji
Hx74EMT0SwrXsjPO6Z4nBLvglAXaWijD9eFgtPQ8ERoP3UirL4SklcbGtpBB7cPEyxX/A7uhTeyr
dBHWLjXhmBpZdB0EddHbc4QKRKitEsOIIO+q1S7U/VUYI6pO3ZF/XSVmjGuzGK1Vy0Fwu0W2r6eJ
xIb6aQAjig6E+IBiRSvaJrXGurPOQpCEXqahf99FedRrK3Pa6ZN8YNMGq6rSBBW9dw6eXNNiOLlM
vMdAN/zFCb9iDg8RKMS2cKbVCHHHn48DDhcyXmBS3UwqLt3AQPVyKo6IUYkdK5cgXWSBRdVFfHV3
41+VfIQDxuI8YbQYvDhINQt+j3Tw+vhGxaec9v2qmHUHl1ZleyI1CjvewLjrn9AJaESeyNde3ShT
LRaZB06Lu/ARclVV2KZ5OC5WiOxgdAOTXmNfnsZXUNPjT11vxWv7lPVZ6WSPhyuuXbK9Sa69v4K3
ysrV/HXW7DXBIYYYKWOVV4Tp/qx63x1n+JCVRDhNKctxPre4J3Gt6OKSf/IoCkp+YMAl58ZJjNo7
E7B+GS0NJ7eoMVUXuJkPZcb9sZfp6wsRWFD67G2u75PL0dDSL69fAyjzQvUjwDiTLx8L+PEjddrh
dJfFwuWGsJpUi7kV/N5u+1VGPkkpodttTr0wuO78CIUg61aLua6t+0dkaXr37k2Ss/X0faWPifDs
xXeRFkD+S5YESJx8mOVpUJW5unK9ZQPNjEDN7gXFB/4OjaAM+/R61yoeJsGGQoItsGqm936y+1I4
cJ/yPWa4KHRFuwqa+uiF8i6QGHuEwe78NVPpipVr/v2auF2mQV+cLdADC0U5JJY1k5mqnxLfNJ4+
dH3LxM5f44YR3gbvOFeCOTgT6pgjDuk8loHKzFVonhbgSBJYHVBZHARWUKKdpxP5Dp2BLns65fkL
dM7IeG1B55TigZMyWM3FFwH0e8wkdQWCpHrC+1gLm+oyR84e0NZU1dir0+rBI3MnKTS1mR45mTkG
Y//qcR+a3BJ22HCUnWBGc3wXJAbyM9e6SIPsyYqXC7+lkQIXSui8szAaqQFO9Ko5ADSSoNDoZSSm
3+MOPY9dNCvLDtXYjFoTgD3z+rODv2CHa3wabEMPDKEEyA2JB4bLB6LPziQo3QTKQcXPvoVpTwwY
HmW2HSpTEqYM4F5bYWL+MTkWK5R0VKEaVFhTTvPISxXnS1IBIu7+bdw6Xq1QAbHU90kKYs8YE0NP
hz71xDL3pv1A45mMdyJatxO0p4M1GmYezfbZ+wRDrx73IFPDfMaJNoWTdIoJNoYU9jl/9qDQNpCr
SRGwGSVztZCCiBQhHpX1rMlgfeFRQT/Zngk7ZIBYgXZHxcCgm0Bts8OGfoL7resiJpnOpI1akGg/
GFobj34cQFbZGS7rcopUa5qV+1SdLqCoYBrv7zPaHwajN4W4nWU5rM87BRwqA73ezJ6dY/WjWoqO
5AmAkiumuezYHMmu3SybMjIhsfU42zl3mjaB8Mxg4YOClqJUmWYc0XJ68PCgJHY4ds8IId3X/NZj
qBzpM9kOsWjqICnVuotx6Ecxf4jjDwVzmzh4KQMz+TVkySGgArUnrHBtbUbIz8HxOBPSyPmvdFb/
N6u0zsep59e6U0hMQzv5dj2ZMzLzjxivKnNpQJfgyruFgR7cnjKgg7XWzXCCIrL0JL/QLfaCryC9
wXmO9jJ8fsbO7AtqEt4NQBSmNoUrtdJGHeR0Un5jOLuL6UPetEZaBj5vMe7z/LPEcFPT4g0KNHE/
/d9acq6srQJtanRtVH7I9IF6DaWJvPboRIPskTsZTHQzDKge2dd7X470IkmFd4GhD8d058O9MtaF
SANBqUDNJ4P6hfEcRoMmJr/wNDzuoYqxZz0ZbaZYklR8/JLoiTQQoO4zsz3uHSAyQdyV3oMEO3Uk
YdT7nPA13hl1qohXooElGsl/Cia9dgE2ucpt/QcyWGoGqt4+CxDXboylkA5CHgIdY1N/UESVijA9
2pzV/mRf8fbWXt+k1ZrYqKBb8T5+pVoAdcp1kI6GYy/dDxMJYIKf0BA6P2Xrm8mmtK9zOX+2sMuO
OsronWf2Bx0bsFZtPQrboPjMqW3AzxRDcMw/yJ4O+5jdGJ+5Eflgk+fd/pir6VOGeRLPBQ/9uzBs
zzANvMtU2beC7HN7hlxz7uxfi0yvZYYlSgmnBsb81M4stlPjByTGShWr05QAUnJ/vnJfz7Yi1SYE
vZ/7ixaGfJurg+dcY50ESZ1N3hmjspsddFLmfLoZat5GuV0HPRUumO0yzRwTqD6d4msJscKjOjoy
NOmnC/Iev0CHl0oxGMFeSOKN6KIB59HOdQC8UsAEyFvhFp1+EU74By93yeYaMN/pisDGHWWJ7C2i
iYtWuP6T5qgCZeTVsNOPoL9mRAITgknla2koGmGz0da2OU4XImsT2CPo94MarUBoQC0eiKrTsWYj
oU/BNDAdfXrUqaJ3zHxc7aJ+D2a0VCeAIJKHNMzP1EdqvPgHagy1lksCxXNvuHmyBah8x+XQH8eD
o1m+fYR7IY4Ss3pLlnQv25Q9gulksr5H/jQH01whLNFpBeQ+vPo345+qOG2Kauf6e7I9ot84O+Xy
Koqfj9A1xfhHleInIVlWS5FKIfdgiTCoCrLBSP6pKixLDuO5CeAnDx8QhjhIkpLQ5mdGeW3KrkYu
a/ZWjdIJ/GrNalLqN6QtXpjNjoe0d2cbwtE0hyY1pHBHnWlqgO1PvoATGffVx94YDU1jbmayAzyF
nkZ/WTyHcCXEDAkSANzLNZWM8ck0nsVDYvvcm+HpW7eKghS8QxAjLXWWSWV1umYHgi8W21UGRIRs
b847ffE+wNFBCz45Ey+oO9/2vA/OaS1ehSuayjOaRBnPVx9hYsl6n8PUdue0Q5IGpz1FNFJTk0EZ
kyCm1i2cmF6pubMtWcGT7wiQ8dsFlhe1Ad1FuzPPYHuI03jF/54Ha0q/iCjTXA3Q6Z9Pnr0kv/Yk
PD4epnRwxGcv2lIa5YYHawQJ5lm18g8Vl2wvqq61508nM8BgHnqMQAqwLE9GYl4uBHbc4uqc8Jn1
lYK5QQ+ml9IyoI4g7KpLxZwF6mptSRjZuWvB4cArk3MPYVHcconQ/9DXIggTCqGw7/lcTSGTpAzz
RXFBjmEucMWq8F5nfMaCnA3+/LLumhnB+p2xmN1jkXKQ4r1JA0W4831E9VGFcrE4+IT/0Rz7fPJp
L4dCzHgABj5iP+HXakeZudkRwZB2VIERGrF3UgNCJs2FLVdgpulDmUxqzl+0xuAhd11RipDO8oJn
LEqtDER2gR2q/8zV8QLjZYH2lXYv+aTsR6ukKcC78xQsYmHhUAgTIB4WP2UgZUNi5dNU2Cs4q0W1
2ectq0pAL9sGaZPJ5WE6h0MSNA9FSOkwd3SLYUaU/4yWhAczu2knDCM1IlOHYAS0yBItA7SCta6P
IVtvX8YCEzlRaDkNm3W3DrPyK9IZhe9bElBWM/TBBLTTdxeuy+5ec7DUD+3TRbGwv5d4HHeEn3al
+9clSbCbm0xcnUz5+K7emgZwDotHUZxRW36KjKyI8cxGpVakxe4h0286GtlISuM33CzyitJ0e7qY
awvLfbgNcYiqY0MB7iSZBKBIBn8yY55F5RwVYz56rZjHTksNxxP2jfBbx4OEHnZQjK0OpewK9Ift
mMdLskwpE01EcA70YTVXVoPTG/2SMdkfapU4aMX2hamwpIqUfrYVSyrvyCM/Pu31qcaThucop4uy
pMStRTx7Bks+TP+BzIjrARkYZDoDeYmIXAMucrVEsRUeEtcTl7arDQEcSb7efcVvkAgbnnpECLDv
F0B5s3XoPNXJa4gmDAjjYx7vJNGevba3APOtwyzIrzIVX7mXC6atET3VtQOEsdZTSgDU3NKo2NFM
r9TxrDyapjjjtKOMKZ3mhjWqhKHxKS/sYvqqemfTsovdyGSynwppHDh/2yRB3x2oEvAjLTi/nJRj
f5H/+jxMwoKI7/Q8tHYzOAJ+QnVMm9Sl21XSr3Cw29a3FqfdHrhV+MSRKgo6rgPDtR2KYj4hhJhs
lyfdVnZ8fVKbRJpOl4j2a6/DaXAhdoRByfv4yS2MgMeffGF7VNOLCYcUwDdbSnQmoTX/h8BK2QKC
QNZaff81x00FB3uu7ED8VqKM09Y4UiZo1RfMeTqC+HmeDaWuWsRVHAX7JskUblIKdQkpT9Trr6Tk
X5FG7wSqUgiSn8hF+h0T3+KTLLJXk4tjzATT/30BSYEwXe/3ZpJaJQ7g1ZxrX9KHg82pTZmrC+u5
+IxstwaZ5r+f0vvlfDrktm93mZWxDwuLz4KrDydjSqWj1IBNKKak1jm34Q3/VvXVzcqXRsR+1zwd
lPgmj++euVs8prX/p844px2iEu28RYuTTIQGdRUvdGxL/WG9TygnA4KCDdZUUkjTtx5T5ZDsbGxB
gQUiixEHNnkgFWIULYoboof+ElgsbKVSH5H+z6lxUU3Lb4kX5uPooV7B4MH6wdTkOTMIM955YLer
kfePkGiQk9sdHCtmnKqrtwHyOrQQz5jAzM8sicoOXuMAsmoRiaE/u24t+7RkKZYyxO8MAlq3XaSa
own1mqWj8FkDo77305DEkLU/uPLyTAxAKeOl/omLwSU8wePyghAlkKrKAc/UR9+vpRad4bRdBrwt
mSUCeo8A0QnbMEQRuEKrmxKhbCshYK+0fhl32k+dQYAs9dhPTTJYRGqqyG9B5xXNlGxAF0gN+2jG
FIn4FeV2T3zyRSGs7jODGC8ePSePh4JTzZvMop2Iu0D0tDMdoXfx08HlwJwmIab0i3wgoBsJfRC/
mjGFRJwMi/lkVFDSS+XrkJaD+Dv982XxB7RXfe2zHzuHov1eoxAjm4kWy2+/mcF5Ksiynh9MXCRt
i+j7lYL9s7gjgGOg0CQdClK6arCCI5Gr2LNqrscKzdXl6hCL9z6B1uGwTFhG36OZFaycvvV30wTV
4hGr86+cn2QxM9vYLiYSB9+I1SWlaMbZIAlYFQEMhlMGpFYzMuZ5zsqEOOuy5FRy+aCQw+IMXF9y
jwq/atNE7PRbPF6yS5k++gOU3bjjsAqXerpfQ9W+hKTvubtzTDFLsJEThRsxqZfuwywtfNJ+o10E
HTnM26Jx2adCixWRYq8OrUOj/DURQXYDklmF9gPCNT11LCshYTE/RdgRFEpr28EJcPt3om0rMzqX
uJE+xc87ojaR08V+R69hkI2fkQ9q6sUgOFyy7DnInCD28Kslk7zwCigSkR3TPDdNleoxwRp9hfqE
nSoIplie7kPyEftFOqtsCNf6nfhJ2d8pRAOA3sHROgWGG7OczPug15/JvKQMmIUJ6aRaHHlSIEGh
XXuRFgbF67HbAa7gYSploedt2LN4nVKMECUVbL4R4P1g6sraXZkWW5JNm6JBVaRUPZi9Rpy1kkiO
eKBUmcBVRjBG2AdfOuQfeyNaWiW6TSDd7aE8nb9QKSRwwurpKxTER+OCdJdiCDF4VdwXCSzp1a7R
vwibNtjgErgYN3fg985WkKM2JPP+NJkZV1sFSwq0E2ZkdxKMwAHR1ZXgcXl6Fucv5HS/dHbnKbpp
UBZyA+2qEJKStg1ZMX+Nk9VVhvD9tfy/SbgOlA4kb8Pn+xJcao9+rwwA8UwmhYdBX4FK5dWJO86g
6+RqIdBPW5TRDGVd0juqxJ1auooMn9k+yynwxfJbmnco90/S/WB4/0AZlyIPkcl7OXb4AH53stLH
i+gtGHJx/gPsehO75WBLMNGUme0w5fJxQKDEP0He/Drs973r0ZNZ71/wokElWHpV+1/p0Gu/i4ml
5nUzIdbSznzIu7GATJpmjRUaDDO/+Ss8vrcvrG+MgMAFAbzIBoum+ewS4mE7Xelg/JHjGx8KlgwE
sQ5saLm1WHpdqmPEmsD2SfAHRxoQjSnu2KkDcp9DReKTOrdi7R/UWDcN8gctcQzmASKhQzwKIf23
wBq/yXf+kVvv0ADag8J+UOsVj2oM2KjPrdWP2xbw6eA9B4Vvic5oK2z1qBlQ4RoGws7Efy3uMg7c
0R9153KYne++uJS4Eb9rxfoJxujbDtcV8YWDmm0O3UpX4cJIuYs7U/49ri39wLZphw5wwDlNKNqL
WJIQ6nKC12bt2s0wvKYWtSlKdtJPZncIgJHeKhy3NKoLVVXiBOIOyfQ2yD2WjnopRoAU/GRrhC33
Tx7QAeoutxhiQygxDk4vBuobrQMbRJaEwCc8yfjOeD/Otmwau2iHxMJ+/tckixtoQfLNgVHQcDm5
/xXgcPdS2b/xRzpUbUSWQG9qY9hLyHEhsG/bl54Cpgjo89v6hvRTrXRzC6uoHi7g+8mQAntr7rVU
59ro2Xgug9QBbDHBMF+UxSGd4fZ+ikT2CmZkIYJ/i509dCyLDsfSnWbKUixZAHQM8jlrXGbkz3IV
PY/tmdyQaWX7nAlqoAeh666jSCXdip5emblbuNicXdcgx2gSJrt2Byo14K+qqN5wvUQ3uGDJHKj3
3pnIV5JDoTVpz0NYb4Xh97T/Y+Cz4W6oJ3SSjrh2lyy1MjJJHLmG+U64lIarcIk3bZ89x3nwn1dQ
7GaMF+X1Dwcf8xfU6WR6Tm6Mjx6HIMN2LhPQ9tQinRP3HfPnsi1ABENm7sOGEqFZ8MQucRbXp+jS
wU6h8f18oA/mmbILTwtY/yllMi4G4lcdU79A9EodD8oKdyvWpEy44r7P01fktGRaGGwySR4ddw+A
xvlpj5h3Vzv64jPP4c7AK5KZeknvPTWFgimNBxqK1Sm1t901E5kV3w1jvMTGNvameJjE67BghrQj
7vDCZS8ObrNaq6OENTypnDpOwwY9lI0yVpy3adCNlsaVVsQVaxOvZJvxV0dhQKmMO4fua5rVuhlB
6LVehExL8k/wgjLrmiXUGEG5XtYKU/wdKXVH3rKxdsLRy4wbj0LsrwgB8cwpvGAVkrkpYgFFd4Gb
R6G84uysqal2qN0POpjuzNYj/b6O1BeIHCay1Ytxd9P0WtknlxLslccvjnFq7g1PQhwM3rJsxBft
y2mP6xnNwm4YTQALy4OK5hXySsIh64MOYWStK6oyFZHHSbbRf0+tp7Ugxil0xEbfV5b3AuWp3wlS
Bv1sncZTlhSaYtDfle80odWm5FQD2BIyYKoLge6RPhpAt4Pg5ZZBgv9Yi5rm90Bghu3OmWSY5KCn
e7qx1Zx4mbUtUyJwuLVa3EpUT8EhkijTYs0YFRoLis5NWIEFNbhh3nE9N1i15CLNhrVYq7gD4yz5
XlTCnH40W2MObVRhwgey8cmuD8Y6eXT/ELPyKYBfICr+1phb+6cK2LnBc1w6ugW6/aMvq8qm2i7F
EB7B6EICUfo6pvhn+MJV7TmaY2WkC8qxjGqUbYUuNsVTqF36yxCw99V0JfJ9k+5X/0lJYM7pGJXN
+b6Mz5egRPERhibyoBpjdkWoZj0J/T4HH0cp4f6ZgErKoPTIqjcqPnEFz8LKQncV33Ebe9SQmf7J
CqNp6nq20/DCq+Czsm0SJVMK+pcam69mhBZhcwjZBCEAEhyLZWsqSYLBtmvJmwAxZeFVdx7kE1Ll
36//dCtH95v/hkwetrboxg7XqoEFQZL3ljTBzTrIWVd87JlesGlb7XgW9bUSgpv1p/ZT7r82AXnO
wwkeeXGxSPF5FxhfYtARVk8cacbjv8IAicA2uVa3J6WCOjG6hqBe3/kk8LSCSVHA3srmlad1Lbry
w7zV9G5y9tq68s2bg0py0ProwO/br58nbj1T7+jU7K5MbXqQJu3OnCwuzH6SrU8kvFsVgnddAP1b
4bwG5Cp9ewhVPVR8GXDi22WisRoeF/+6xzN1redSnBpRfVqhhepP9SL7jvOb7O7OGE7IFHzrTI16
AFrSn/eBfyOJw//YnQFPppDuB6/iPgBpiV86mU43hBe/yFbUmpBZJtM2hSm+pIv7SYByS4sZAdJ5
ubzCfh41APXc8TwCJl1j/Ja6BDPavMfMD7SRzaHZmOaodt+8MfmFJ6gTplPVL8X/v8EJmH4fPLAj
z7yfprE/brDa3hqhmYmOD+f8xG03Guy4DQkFVwWOinkjH7J7PaycikPN0Y4Ng3O7ANHw8MjCl1hT
IYDIl32TyYJB3xc+nJ08eSL55YP0ExCOBjPlXYrRqPVjlr3Gn+yRaatgGsQHa567Vw7epHXCUZz9
A+Ikji+L+MjGYnoXL7oA/VLbuxfSj3LW//ZHenOGENJZG25E+OWV8Loy6ZCuKMbV5DkpRoFDEHwj
oGmT7nfjHtUd+V+rO6Mg6OAVp/HDa7Drbwr9AS9P317k8XLDEMlJqhEdEy1RPVnANWOc2oC1W0rU
PmwxeVUgId8axoiUIsg7r5Cjp05aLfAOseC+VzfmDjBS2bs6KXODbNDMUz4Mjiy8cFE6mopb/Exm
cWaJyko/nhNkO2czvPYkL/wbouFk4P+F4qtbzy02GhQnFWBSN+dxn8z4BgYZdOVcZYhk2JB2HvHf
KWCHCQX30K9wmOLsaHkhDC3CrN0326oiIoEdc0AhXYnoWH+NFBvxJTrNoPxQPaH/++Vze6Xvx2L6
SRN5TJtfnr/ClcDVaih/rbfdkJid7GbOopceJgAvaTSO86MO1aXd+H+Hjq6se2txY8N25/Fj//oh
4kibt4k5ydoTGvndLIyUVkqfD/UYXwS90/jPpbQKkiVc6tWSOX6aPEeyChqG+fqeUM4n+TxkUKfj
Mx0YdkwXKaY/xmdguZ1+wCvZG+3sJxoRaYw9BTFj0nQro4LDkALAQX1ZagH9+/UHKYfZ4BBG/IfB
NDDc97u/WIED3zuOCZGSSDtnBzpa3AD3tyZKkz4RPyEbSNKiwM8RIy+20HYQ6GJK8/T5yOr787lO
exxyGH8meQe+XANsBAfAevRYRmg3b85fZGokO5wkDNR+ZGxWli+aXuo0K7acGZQHOWzufvYumVYV
173/K4ldTwMPPlnQYzqnFOcqn4NfhmpuKywOZ41JXNimxfDmPi/mZkzzMYVu6ii+rsTsqCWxSrOY
/kALgltoWM+euVuS0vH3fq6vAiDorHhCJxdR8O/X62ndJ+p97B4NfG08/DwfRoRLJ2jjdkncG9uO
WS94VNGp9rL90Ey4EoBG7s5sVrJW/xsNQh2lK+CnnnpjcvTWDruGsz0lrX0J3RA2HgzgDZEq/g2G
M4l6Yqs+C8i5RM8At2Rs7Gsd0ykR5jDtr0d4Bu3G1nqvGnlrt2hU1xr/Xpiv7L7bwUy92nFSzkjM
srbL3Jf8VFYctC0mpgSJwQ7W/e5Yvn6Nm+NF5uoMgQROwTCk/9kNpIM5rGH3b3srIDITU+ld7MVj
bXWlGXDMEPs0ioKZiIsYvTbKcUSlsQdLQyaWFDgo8FngVzDDQdekpO/Oj/LrUfsbVtbJd+cwy4aQ
kIp/Xg2MefrSqlPZ4SReDjAD+LNdX+JCr3Km90hSahRRMEiIy40HXb0Y3H4Sw7eg8mKlUX3Q2a2L
yoqi5ubezWr1KA2ilRBrZWPqYCw9chN/mZnQvitPlYh5HE6VP8Tpk+LUcC9baIP/fLDWGV6orxph
YCzLpLGiZIISwMewDHz//gy3V2+Nhs27WfcdGB4o5ghkOR7BHd+gjs8UytRyv/SSk8hJryJ//2Tw
OwUOIHgcaRwt28Lqm2FlWajQcjrF6qieiji0rcTrGvCKmC3QUcjNorBZG1Nh+NljyURXkp+u51NL
YKn3vQ4UZYbMAr1XFQ9tDqjqMfL4KtbxoQlW+uqSkeJgf1f1U8UwCl/RS7VbM8CiwFm4T4B7Y9fL
c+RkWBPczEWV1me9n3oBuv123Y8MxLJ0A9XpueIeoAGKmYeoHaJ9cmxwi4TJge+XeMb6Z8Jirhpy
GyPtu3fPU6ttKLVtwOLSXRl/EsShj92FytaZnlbFpN98/GKQQGqkIWDrA/N3MGyZN0N88ei4hky4
bKM14CCeBJgiGvPedx6HcLCAnxB1EUbn0UcmSP7pkaPBEmSRsL3deGFS0JhKMA7kdYQwM2U2Ug5q
W087lDttMy+OHx7MabUBxW1Y9ian912speeXbs5y4Tf9pRrCpLyilSwhzWTevZtCXO1krcXiv8G4
vbCowb3W7vc7VblkAwLy2R39rhLqfqf4odYBD5fLIL5CHTycPLamS4jD7rw/UN73dQ0PmpxYabQi
U1fq8VFqRKYrMN819k0dEvkFfPFHW97WnitAhze5uoV+/vinSLQTesjgNiMn/sn5pIAU6JUwv7gx
hcoXp9XMeFVVnSDFyCrYoOguY0hFbkdNgeNYZdTaWP8su3NJ8uk6iLscWyob4wlAkUOnWT1IvIO7
OdcyZc6rwm/ettvSB9Fk5R5P0ClVjC0U0DIsN2DpxFt9cs41utL0EtLe44CGgacBXJ7JbPOeFN1i
9QRxme6IBz2f1J2jpJG6g4qzPpS/rZ6wGkUGaO48l8O/ZpdHztvU09kDOG+82imDQuatQSsvhqRB
YPcMDZm702AWmV1E+l/hUnryb/W1C2eilgOcq1fc7aPn5k7XOhR3NWrG4aUp+01I5fkWpi3A9uBk
oHh7XYy3kaqm1ZAoE2/GyIUN8jCFY8stXhNOwXj7ZQZ/AkmxMAAGpgAN5CLxrJuoRUsUg/Ety+l4
eJ4cO45ZeCVdXUlldDR9gQgnqJdpHAEKmWmkdGIMlFjmfouXKGnq/q91Ir8bdqwu6E+OumsvUbfK
NjxnvmrURn/g12kqYMw7qWaXXAY5tDZoXfIUCPZowPF8BnXOUkocJJHOukq3tRRVFAC50B+j/Fn3
vCE6KnViHGmgDpckKnkCE8aaPfYDl5Adddl01BG5OR1plgUEVWnLzMXxqEcFy2EyhFDtbVeHonuF
DU6KWRz5h8vM9ds1eOLVrXDcv63UxtfUhgQ8GXX33IZV13oRqQ0NC/55OS0laMTQB9l4VCKIE4jK
x5p6q0ncn4GOWyZy1KTbF81nu/qOQUwlviJLKw8DcHwcsLNvImxZvR+ykX77Hk938N/NZme6YBHw
TqTHhGqdIEq8CarwbexE54Z/YYN/Ro2ncanPjtuBwqQIK/6lq0+OAjwrT1gEMILA+quPzv0oz+pw
Lqe8zeXLB1UH+6lYEuBQ1ywvWj4DkOIpt+aymAQb0CQln7HTTzR/5CyRO+X7mc4SoP+FnWtJjZKm
L6Rk4yd8972ByGoRrVcrGFjYp/a3SB4JxOK8f9VB96XmMVnkq20C318Og62lf6BwdSopN8tiBcSx
5GFTQxePuZhfsU2PbTGvV+wHkXK0f9xi42GwhTKJXCFfIPrkaed3AGfiqZnJWmmxuULxK+E29ApR
/SNUiYvDv5jbmcQsRt4StgOqibXyi0poDY/3uwsZv+3iSSGVkWTMXAe9+0su8hHqb2sU2AIXHIYh
oZ6hM1Qkg+4BQ+w+4vfkupvJYEjGNtfh+3ibfbDj3AvBiK/BLS13Xs/J1nkK4xPZaOi4Px7LqdXV
1h6KJ+iV2HuYhwIMTfvUP7MmyhwTttphROyMxJ6FBQqbh0dRDdGYaJsV0iFjgPjmca+ggOuRR70d
SA4GeltZL2m1S4DyIjswT5bMQYRQqhpGUw82wGOF4UP3yxY1P0cIsYHiOgdKugHqTgF0qHj1VoJy
Zux78DqY3LckWPAJDJE1++/4OgGcDVu+iz7gKvaT1Bmia37+8Rhgn4uAe7FAPUap1qX+71nmNaS1
hXYIWLYmAgYgKvMaolcaeBvbvKs+ZS/ja1fVHU8yKQURfC/KOhbA2Y1JS0A0WW0pOALlbQRDqxbW
btvv3Q8rzXLs/jV8d7dc7elp+6cAnRT9/G23kI93RPBRs0a7bKXAEdYYwsjfn2vHhEHanGX+l1AK
X4H1rAwHpiPvxFV7H8PYXe63CHMnEs2Z+AwnOODy80cY6lkfplEbYQUr7fYVKaP/f2LOn9Kcrllk
ZSMXWxAig5S4qKdfWlaE7ZN9XVnp1wLQ9e5xewg829q7u/Ofi4d/eOLjPqqbHABEYNXQ1xvvpF+x
e59jbkoqZqla7oWPh5Bx6dCvx4cvxAF4sR+GUYSFOGVFEnE8B7vLjbA6Q7geHbargBGDH7zo70yG
v+OpX+XVMWmKkg+7LVI9d++uT2TionNlHpQp6eEClaCcZYvTlF1LZgGuKA9NvPE2m1CYw4QU3yMq
6BtfWdpNeLxghW/HF59tUInUct4UpwCbgh1TcSTeHyunHhdvQKY9mLvp24C6+VsZ1hjpGdUiDJgP
Ll15nusg8CNhihQdR9Ykje9ZcUXQtTHEUzERwcckZ4AofKbwSKRd1ddHUSitvUAd/q0T66rhsMmd
hAaWcA/+UfjLf9NYOtuRTsxZgOt/YoryiIGfZ53AkGJrW9dG8Dbgzx9eQWMltz75sb2x0ohueKmS
4vPGm03GRG7f7nZj0og/1YxgREIqMIC7K6mlAO/iMhhn7RkFFpl8+cHmx9NSwHVvBmHmquqSLGLu
5rLf+1zb9VhbMJtTkNJAZtvn5Nyy0ncpvPY6LQTo7N6ypu3jOVTCFJ56sFiHgiQJr5Pfx1h0GEp0
2mrgaNrkRzOh3Ybjxn/N3MygaiL1JOxEDIK7PB2IORLK0HkBE1v4FLBGC9M8F0fZv0C4lBzGsL51
vYzkCqaLvkH9WRQXmNKlGdfAgkieBPikeCTMgcHNilBW/NsaEu9WSIXgISH/HLrFdXfaIvOaO2kR
5JFJgnHYISHj3RBDqSA19K011Dgbcy8LSpm8cdKces71Ktzh/oiDI1pOQlfM2WDnwEN0nesYUPQ0
Wh4ZIyL0TtS7I9jmfq9jFoe/CHZzJWaHFci7C5MSURx894IgBPV/ZhTq4inD5h9e7ey25sZK9Gtf
N7fV/4tTV7ly2lmEAOu3Bf9+T0EKZS5aJvRrOfYGbROR968ZNOvx7oHSsw2zAOjc2bbgVVi4MLb6
IZl0Xcf778noSbjklL0sLfALulqUJIOt8QeOXX+PoGtS5AhmjzWPCerW4WqLxA2l6l2WiBQRzabH
UHGrJvMC3QflAMJ7GzZvXDe51MIbSooEmh0Nu6F7SJLc3e6mW04uUn4VojvaVARMDSr8qWQyTfUD
DXsDVlKcEQV8roXFIcjmIrS7p+8ATUaZv9F6rgkUvIh45YZOxdOc7dkG1E7XwHdZg1z7B0reQgtl
wx0S4Tm5yQ4h4/J75dv8SNG+bH+hiHXjs+ivHTF1h4Pc5rnOIF+erWRteZTGbz4wDM0OHqZ9oJR4
/7qACM8Io+Xog4oCi+jNrUf5n3ZkIK+Mx6wrReMkXTmR+AhIodPBv+eZk9SD36ovbQYXUQqrcARu
qQDpmmUfl8ZrbB3ooJs1D8meIn6HCw1C77m1P+fb0fVoOZqpnUeXeZfpZ41ZghbeUkpfCB4VJbO4
lXg+8GF7RtJdMpK0Gpcj4gZavRwxw/xD5buTqZcRuSYi7VugX8diPrEzWfesYLKnTPr8vDd6Qj3H
WklafuDbM1eB49KvlW49NgfGVYVbt6evN4o93g0XcQFVGWhuPBgOZPNLURUJneN74Lx16zETFU2r
D6+bktI+KWXMBgn8IqIjKPButiD0C9fvloHcsHHCPgsuKQ1dGms21kBtwJFptGmEgzpbDj10TuyF
tFKh/NI+WXeM6TVyUGvdQgjD7oZzFakcAQ13N2DwFVMF1eQu6Z2Cu6Jafo+Eei4+aQcRV+5y9cLq
2zBpE+2TDbh4MkdhHFw3aYvu048ueCVQNvZdXIYieHyJf3lhCmvV2+IaGuDkpAbmNXnOgiZruY+t
9gGn1FtoY22AtsiPS4SjTgz0xMFhvi6LwFz/zbQC3JEGLxJ0VVXmHQhw0XdDwZsOlytYU5LLYGZn
viTvs+ZeVemu0aeKAp18Tq21tvyPCbcGVYDrlBh14vg6aD+9pGtUeZsSOAD6yIX9k/tvaFxVmxum
65rzATJV8iXHgmbPXwFa1sf3MsX5Y/PCdHEOd72eKUCbGdQgp/zfXtN5uD9nkKCxWpaeuatoEvAw
IS0EPuGXAtfXtR1j/evW9kM8Dl0OkWuHcRWkNMyDT99G+sYrRTkY2zk77g8kON2I4lLCtDvryj0r
8wZDJENBZNhv+2L/MeCDJACaVx4VmkkeqhmfS2WGAvumHieTfPFB13NtFZn7AlKwRLaUhSx3MtPd
/jWZSnbWM1DejDKesZfU7FpVI1d+W92y8azzVQEvIvEqjmMLznI0oU5idDe38bHeQc0gxQSnh0Gg
MmZPx6j+AopUHfbDw2HlPN1UHo5QDCs/HOUJdqL2WYd9VHfjZYRIDj8KOzDfqBKM3ws+t85eSiRD
7ix9M9OSoaqR5xh0ihLWCK4nXuDpHbaJZE5b+zzvc/2NeD9GEMwOuvU/lZNPajM/tc42+8LJpQFp
Vq17Bl9OTYlXXj3+4rMqQ5IROQhWBZpHf1ciJoXIN/m8Ef4shMuI3om84zkHR4mEGLGn75zfdkWh
nuPmdn7x+1drjit7i1l0/x3XkNB7QBKczVZat7NX2a3Iap+DkM5vq1BziVJ863O6jTl0vXTDh3hh
30HYp+df+VeStJD5ZwQbmiB2s/RVEnIqcTvzOXvk/Q98E0rxXSL+n9m8GS91q6iIx4ywngRpmlqM
y2g+vsOD4eEOtlWRIUuMoj/9zP8hgvLd6ErPfekEtKHd3FyBfC1WxAYLOBlad+twKVCHEZ/6860T
SsQvSKs/kVQJLUIruCnuwaDVh3h91vSQOMLhVDOMJ71jfWFvvF67E6RtDx/mqPbgOrugmQAe17Ge
9mw80JzJHOtvdFvZYAJoGoAKOFhrGJicsTUv/bt4xRcbFOj6csS1EgIGyLoLrSt3o+7GNc+cyT88
4r0K5PyKwGnjVrZWRELvex/WRdjfjCzcF7Oc7H1HEXV8E8CXQySUwF82lyjB5QhGsMMP5a+w54Nr
ovvPVc3fUZB1QKwUsPLfEwgrpesRosrL1qE8G8JmldClEQ1Ok7w0UrL3J0OY12Fuqi4hHLhxUpsz
A7eL9BYIHZF4Z52qU3QLltGyuJBhIJmhd+IjbabpPr/+UryaViUXplyrTgQSx+slIquvkrkpg8aI
QUmwbQpDtmLqyzZhQTnxWHn1o3Kpx2TMNFx+/g1Yo1rfPMvF1GsMe6/CVSod8ec5HfGLIbKh1UrL
35GdeYIoOvutt47oIekpV2GHiwZmX/y6UcdhBifim/yzdPAamMNFhCNJQAPHROZFQXETH1c6rbKW
P5zYUryqLbEuzNrgqdpJqJqbhG6tetYnAmCusc7ImLImY2SDiSG2SJGudemsVCLCX0tibR7ZVr80
UzEKGt6DMV63IL6mJ37Ox2o5aPUgBjK04fyiZDBwaVJ1yxcCHOOoAtniXWBg+5oHehKEbaWISvAz
uz6ysif6CuoKycvd78HVAj92fJdcC/egYnIFURgshHTT9PzsjZkRVskiXHoDzJaSWZt3+7k6KT1Q
0x+0TfUmO4kL7cFNk5ulSu+OS8+4lJi+wpuk9pxsNDSYSUqF1TAJehmj/1xl1UCHRXLi4LW/QyBx
/n2HCEnYF7pJXqeM955UYAyYeNQ+iNARpUZwLWjSfAnLIJRc/CesLuT1QAxmixZ8nkPSwsAxbg64
kVCTbpOXZfmoshuGoYam4kKSFLdP5ZhtmtdD7kIePp4c8S4e76rTxLBVZScBBLFmJzD/dg9qrbAD
40KFH8JF/rLcZg320Qwwo0lXe3rkUh0U07fpGMpVZ1WuDp1orpjTV66sUS5GkOt87FkufBL7IcqK
9MsWVFMkQtXQFHaC3dqV2vrckXY13QxxFAonzYkcMVthawCIphVbsOOsAwbBNirPaK+Q2i3wHLFm
kP0Jkc7PxHD+SwGgoUuvcKveQMBwqWaNCln8OsWOUuuWF9LLe9OEqRKcMDT8ERQg5NKqQyxfw48d
Yt7EM1aIHHEzQEMkmXywkvLIZ+hKZJRbpRR23pA3go59nwBI/0jZ0NRr5qznPxpJ3zjL6PjP1mCL
lr7JQRmul8AKsQsGFd+d1A/BUn9fP6SMkEVpXLrKW4wOdoAcbbLvlmOnhqOEP3S60l/Sd1s4IJH1
pgHQyB0vdPIEmj705WIE/tZBXcjUFyp2Ryxb9kBySffGpWdquhHW3D/Rjie8Af7eLSfN8nDgLU7v
OgH39EX+lKZMQ6dCkkbTu9EXYI0YATzgW0MVoknmhG8Z2fST/zr3pPz/85CGqZul5oimqacEcOTs
xaSQeuY0s15MnJHX49JmM15dWFly0yxKahZizmecBXASsBkLMXkMCX2RpTXwUA+awgut623cL3Ft
aZxuSSDmS5w2UqxAxiv5xVIqqCuaq4h2s416f1nwYTOYoSt5yAu4tc6qk5Awy+EbHlN5kDZZAeGn
OJEdlZeXICF8D5tGHf6iLz7GAizv13pk5Z01xZI0V+jn/oOAZxoCeORGcb+QL3u564vEjGl9w8eR
glCXFQFhbrrsVL0Ns6wNbrfpVAJ05cuciiac+FjfQBZCkzBft4039bMTNHr7rXhBIuqE93XRXrVa
viHnKkl7ce/+PrP5fXu1DFyCbcAOMBUPO65FdDldS+y20LypdnN0eK9IoZ+rEE2qQ6TFJIS9O/iN
ADJuHZtjjBEbEL5EDcuQ7FFvAoLYLTnnbHp2BybBI+dBfTaxrK7jtwJbI5Y6BRdswQmpNRz6Tr4J
ueMXXstVCQWFMXaqhohvCYMVA7q1GxFNvInfCxtGuOI5/5hWM37g7FpVbNbP0cTmW3RnQ3PclG63
VhtFE8TbtXco3nsmoG5ThykDKLIITcKqohnaWR2hoKFLPd8cLrlFUNshtWG0OnyA8gm0EZj8Swyo
S5r7qFI76PLiIx90gJgSLrD9Mzsc3hXV6omChoOZPIvMIRVEu67WeAiw4z2goyyRthAlzeRrDFT3
td6dwxvG+GwpJdJxKDhTrF5MLPkiSo8sZU2b6M16HiOyPlish6n3aVQ3ftcmOolaKl732jNhpUhv
5Lk5mQF1OZOxQyPevSS4EtsRSnBSfXe+Er92lRKxBlE7zJmXQBXpeGhGs6ek6rXHt7Hqfdl8ctEP
TO/vVmEAJlISf+SyR4zHBDRqoWfYq5Jv1domaLw82GJnQd472KJuxkX0jK8u5T8ikV2qZliXLYjA
7jUqDPUA1pGnAdiOfTR5fyclJBrYI483HJk+v6QtnVOaTqIYR3rkNJzPKoNNltE2Uf16Zs5wak32
dQhbFG9jvC+Woc/Pt/dKqS856e0rNg1nQKGS32DWW6VXFlqOnhydh1+LbeqwE5O911z7H7GvyLXi
braX0bQV+kuSivmQTDLVRE6xHIpjfIWhI+vJNKoUH8w+hNA6fvPkKDKxoBeqxFAGhkzjejoenRjl
Z4YIxhUcNUue2Bx+IBLJCgoGAmBYx0CsXsaoju5zC7j1hs1+Z7C85mLf4smP+QFP+aLPp7vQYc9B
tSM6u6UlfnWaS/yfbgyAIjLCGCWmozMy36r0wpBUezRwsMsCJanslh+c25P0jZDV7RKd11HyG3UL
eR900DkPclJ5IdL5SeLtccjmqoXq0eomrznwbULDU+uxe4bgwshmOrITSFJOV3cb9BoKoAqZAaPH
bchCOxeF8qL77P51PyM7KliC5k6tReBXDVrNAtyBkP34zwlE+k2e6hGQm18kS8XOrhldakg3JyCM
5STnS2bVwb3qoMoTTJnFh+9Bj+dv8TCRqNH/cxpZ2gCBrk6AjH/2mqBpylG0+v9cNtbfJMwO0Ui8
slmB8rd86n5H8cZe/xMnVCvNHZn5hC0aBi8dSgZrWzgaKj14xcMGkrz2bCUP5vzh897Wm/iZnkp9
squcXWKRxDdcf/L5XLJ9QEts9DW+6D1dKDv4cTBI64jSar26ztJacCAMQTYoEGX3QumkXyqQlb1V
ty0TbF0xybvNO40hG8N/zC+S10WHPWsMs0xmCANYomexkQNaTovUxuxt5EKscc0J5rMtu39/MJl7
c078Oc29NVdwtnAk7m+vzuu2dKHtxpJuJI+H6TCJ7OQQU1zkmP1wVGyF1GeWXjBip3R30uTnUbvG
w3+OY9ZgpjY7M8/NnjtlCCPjkQ28eBeuwO73VrwI3c4uh/odhgFoLn5z9bfyvFspYXBD3wltbkOG
pjZPkh8S3pO4n/p3nZqoDE7K2djYEBtVJUtLemDvBxCgg9ItDOivw2hnSk0KMqVdMjlwoSuz8L/j
Ik6xvVOEK3uD5eA83fkEMu5akrI5dBrQeUCqVPW9xVIz605XeTsVz0317NZ0GcDXIqNWVVw4uyQl
jolp3AmmDgPhcJTe60ErkKIF9qGmS1fXqFE4j+xmlkwO6IQ3QtrkVZ15jV0q3OftsN64wJ6F4Biu
Uqko3vvbxi/+ul/YbHoyITBw8f6fp3lE7gAvHbgqUJjD0fJvA+HwLXcji1RXKqtARI/oKkobMkAy
Yrgl88aFcoWQNFDVcfK+wGBU5ZAJiRfLvuR+wGy9qcvJfNI9ewW8/EIE/be9QdcT+dp+cRzmCdsA
0ngc/XVGqyu9Qm3QMzfQ3clQn5yJCJTTlBxF90ATsXIdrcNmdBEvwHR1yEoSU8poOHI4UE/vYgU6
uW0NtCwMKgg/EWUOzmP4SLZNSmqPae8rwtM9KgFqkYeTEg1V1qt2kI8+PBIZQ7ZhIGIryCaDGlMe
3z2eM5Xw5fhjKMCH516NUNVpr5zV3cssgpXH5/tZ9C8GgXE12lQNyzbcKzlfaR38mZHQyyG/l1pF
cLdAGKgVyo9IF5I3658HtWZleM7ONtGdIb8cOIxh44VCY/dySa0ekDpx83cVEgGmVgvA07n+QU4H
87IEgQj7C+bYCKJWgv328HoI/DD9gqYfxv7mp4Nscdo7+f1+b0WBj34MtWJ6VRnbHepsM9MuefC0
pZk4EQ3Q6PIPaqzrwObou/pqpxFi1+MJGUEh0035waaR4VFNQgwcNo/h6+QuakIRv/HifY/qPn8A
Yy+VNZY2si6E3Bis5oG4vNp6RcTViQVw2dwovuUqr/TfGgBEFSirS4Wxrlm0WzZlpVIRduGySCqb
gxrcZNNOXUCMtHTkbsOj1YEObR+I2t+dNZnCiDEd1VPzDH6uTZKm66Nm7av/zP3L1ivQB001fmm0
xmT8dWzhRnquZUsjTwwnOSdiAM/lGqziGXesRA+xwFkA22KJtALM+VDIFZl9AmILjeSeHAPkl2LF
Xfizh5Y3DaUlCG1r+LrNsAHtMKWqMGQ+MQcOX1BBFsRcvskRb/MamEd7ilfcFCEeUroXmD6QcltZ
jDGzW5RxacZHfOgivuunU2mIzxHRYGeHV7YgG6/D+XSfp74W71Su6MNsEXso99yxkua3VV8vSjwh
8Pv2UKBeVHGNhB6KCndjbd/9HT4BUxapJupZbhwaLgCdBNJd9hDFrMdWPnxsckjk6VHBPIqxitAb
ceC/WvGljO+98uMCrIc6ZlFlUlPNO8sOiHB5nuRRX22e5GTInQEMLvMZsFGh/DiRPGI1qs18ROvh
E+4bJ69t67eYcTrFfG37Tr2vrOW1iuxE/8jTUsQoJmKxznizr1qcBREvJLHzOi2sj+Lw/DCHYjs2
H+KM6YxwsF9ZX+PpfNg+2mqfWlogUSdgUyvi3IZeqc1bsrDpH2ZiMiZzvZdOncigZ+RLTsu6K8x3
Mah5BuOP5Rt0xgoYdKpxicKHqTM154d12a3igdiiE9jdPdf12UUNyf9rPNpv9ToCvsny9LLfnNUI
tqia5JTrobWLdVV9F1kLWthpgrLmk7/QzM1Pt8oOO4BLkwtRRzF31YMhKD2uouDh5aS+RqHCXnUA
Oo3+iAd7LyyZ+t4geNqEV3zVZucovj8XC070lX2SdFq+PM/bkvd8ZTdRkoEJiHKEBVl6TupCMUMl
KygCDjfuRM8UAOtUrbjb1kyiDd/fb6G6kOfqAgyXs4IuO92F2gZg6bUdU6p25j6wf5+g85ayIfok
Ba+Ort//zIBHl6D3QYIrI6vzeCE6hU2ZtSzelmyimnnOdi/bThtq4FSqizcKMJhsE2pLcO5mfYZ6
cfSNFf9grhoDmo+uFZBQvWR0d4xswcUD1fCGgBBfC99mqZOhUsCOBjJLao2mqHKbwTnMXV8MfXB1
NVAA6vXXpWN83QfDPbXFaHtVKC0A9zk5KeaEgKNz0A8GSbXI16fhBLhPh7VOxCKsz5zHTkn01PDM
zCm+bNNeRwGttFBZZAMUwe+ED0WJrJVyw1c9qYLIZkrppfabzlLKbKucrk6nYYlTQs8qzQkm2MWi
FRiCkMZ3ZGVgG6vjY/j0zM8zOMCbZ1GLmF0HRFOTrVJov+FewV5VWyyAO6m0FG8v6EJlSaq2xDFH
tIz0KQf56SDU8tXxj6ENqDDQ9/k2XhmWmPude3k/6ZWdFJksOQNheMT46S3s+9lWUUW0o5gOzML0
d5psaZ3dEIICqSRuGvS6q4nVv5KiXlynHuHKY1Sx9E8p5ay5MtgqG67LzGxOGtC9iSoD4agrLuOK
f0WNgCJB7IuBLTHrZJxxJXd8iWQDqBBVZUI0P3CEIveV9jtkPgNc7Pnocc1BMWaxAHNRgS5usG79
onuHvM8FdM8lmx4Xvy5bZuvql4yJ0TPPE/EWJBmKuIUcq+6b6ve80DID+e6tGJ5hzBl+VSb8dn/R
NFD+ULzQfv+VwZR5MzbRCOlZmHdAwZzyxAs1qah+5OZkmeC0cGUgxR32kcwwB9gbHSYYys4tqdNu
ZIuMjA0sM9Wt7N7XXWchu00DWE2iiP+KsnSqr4WxJFpQExnXf6E39WWaLjnNq8yUolfVftAsnAAU
hdE0T4Gp0x5is+1t0Px+3ZM9dCVXod26j0MsFncN7twOn4dO6G3qNFVieagNCfOFtSI3AVzTriUy
tSG+7odGzBSzbIJKdMiODGoevMv4JmDq5mxlGg7VaNPpZ4FUsEjIeaVaorTsHiuPYd2y+flBk2As
eh4djra9WvwFNvKhXd+js++rg5//a4Xy0nrqDXimPRPee77AGJEW1XdAf5nHQ+Y3zzLMXRUMDKbl
4sdFlK1MptmeVvCDeZK4rjRaTYpGn1ItZCWsDnyjX9k/Si5aiIOgiNW8HPnE7NG8WstFnFZ+/6HA
Dn2d+peP2scU5rUvDuzqD3T4N3OLJ/5sYdLfpxW16yku8vRNiygclA9eXjgGCmcXjNyqa8rGcCB4
JX366Smg4b+FF4AmpQYtM0PS3AqPiUer2UHfP0tKVoNVppIV/lDumDSd8MsXTqoZKcdjN6A1AjQM
zOsiEw6pk4UbA/3Oxe1PeXdMBZU2YkH0yoyra50pp75PNBk+GfgebCnjiRUBhKwcddT6wU6VyCcz
H2jwqJI2qq5wjljfWRKPYWfciQrAIHcu6QxOyjvKZNhKrr5RBq+uJbG/zlLwYbgLo9XyeARIxsxj
3nzlXWeD8ZIuCWktdS6QFIJhSSpNoArNyuOa/BUfCmJzv9CYksjnZ7ooeKcV6Uzxy97Ty6xS1TW5
JemO/jGQ9UrdF1e9cg6wi7/JWforUV6AYI10LJo5nKfMbDItwYQHB6rSzYp0DtkzHgl/K4IfrAf5
xBaul/7bDz49TLdOm8y8WovnIlFKZeezEnFQXuRCneRfH5dtz3WJbbLtMr6wItSwYkSfjBEXBt9r
umL540SH2hpWMuk1gCwpLTTh6i+C7aZ+XrLiM6reTyOg5La8LU2T0LPm90kwBit5fk1mH4dahJW+
Wx35p+vwj9ceSxP48LIMW4nE5StZ/NNcTYaPZbBe5CZtg0hkST2GwQro+7g3Ph5pCdLHnco/+1CV
YH3Gz1wK6qExIgXpwpHT8Xyzq6JxT36/Id9cnnZ2wrydOh8xlm48Ng==
`pragma protect end_protected
