package rmap_target_read_command_header_initiator_logic_address_pkg is
	
end package rmap_target_read_command_header_initiator_logic_address_pkg;

package body rmap_target_read_command_header_initiator_logic_address_pkg is
	
end package body rmap_target_read_command_header_initiator_logic_address_pkg;
