package rmap_memory_area_nfee_pkg is
	
end package rmap_memory_area_nfee_pkg;

package body rmap_memory_area_nfee_pkg is
	
end package body rmap_memory_area_nfee_pkg;
