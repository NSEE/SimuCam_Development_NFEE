package rmap_target_userp_app_pkg is
	
end package rmap_target_userp_app_pkg;

package body rmap_target_userp_app_pkg is
	
end package body rmap_target_userp_app_pkg;
