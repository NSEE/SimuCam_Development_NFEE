package rmap_target_write_pkg is
	
end package rmap_target_write_pkg;

package body rmap_target_write_pkg is
	
end package body rmap_target_write_pkg;
