// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:54:03 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OymNAx4xY0jKWruucbvRU0PcjvTjCRMtBaEUpEMtl3EBAnJY7QhJ/MNL8VMfgGNe
Vl65JsCUh/rDmk1O5sQZR6NLzGTutJiX2ZRifZ40PBz/4SJ1E4ywUBJLc4mTZd36
IFI4eizgRiQcfWD4wBSLy1VA1XN61B+EXoIYXOn/LAY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5712)
aKj3niifZFYU+YNr3t6aUhVCKt9+6CVDg3ubAcZu6jznenua6CbDP9D+LgCYxZJV
eRfZx/qB/R4P6x+X6m2bvAWlIdydsfEiLotFJAN96s7UYw+MYdFcDChAtoZW2hVn
uMM7qQFYgAypi9EyCk1BE6JGWtbRPrKHtenHXPZjRXmy723HYqVlWLQrNcj2roTE
9K02AkVs6ZBhpTb9M5q1ZOjKbHDbh6IptsNv03PseNZiTTYzYSyU84CT3OOE14aW
M/cH2UNzciG+1JEOfqbPP3Sgjb1iHLNWHSxMy3AD2zdh/8vmKrtr6y3IYCER/gYN
YhxDjfZUYkxC8HMPs7/UKzJqfavjIey1ru9Y1V93xXcW29zcd7JiWiUm/TeavV6G
w2++eQlEZ5LT+KYtyQzBY/DQCXy1hlaHoBpl4btCU9rBhQWGriOYr/XK9cDAmTVw
PYBClm0twhXD5K/SmH6jYtRqYq+sybTgtV08NpvlG4FpcEDL01dJNcqvtK1l8oB7
lW20YccpXgwcz6RGognb4+9Xw6zPiM3PGprYkn07Nm08JtOhnsJZk1sWPkyriXNK
icUtVWpwSvDzuDJNN4bxII32Z8wcSDqb16pOihsvD4Tr0Ru6FJD05JVkK7Vuewok
VM2+RIp6UpMrW4pPUNPPNQDW1v3xVl9B12/EwixootNs6+svDX8KWAY0GJ24ATLR
TsEfFvU4/kbRFd+4bEtX8JJLLHcEosiDCKS4Z6ARXULLrDNqdOrFw1lNVdviwB5v
WPRxfjzyxmvGDu8V1eJi3D365bPkDwMLRnYY9/o/DFMnLsADDCpZQba2p8SSpU6M
Yo4jng63wCNZDOKesKt8Qnj6QeE1csMMXev/H+eOkwhh9FvGd5tXHAohqwQOw0y0
HYt7wnI0SPyYygpiT9NzF3Twy7C30mGhaQbyOEqbYTBESZg5T/cZ0A6/ngRpVxgR
b6zup9CwkJbmpbf4K4xONlwrUvUg9TMzrLjAgAkFNkJbHtsdfksisG9sVruGsZsX
xT5BF8NRJB+1XHJzz5FbK1mQfMcfJZoJ6GJwWxCf0SunNHsTB59eoRhHjnf5dMTC
ha+zx8ImIxD7tePmaOGgmOrUX5myDVwAOAF/0K0CVbO1TeTM1l73S2Sdtc2L4szq
zXeSaP2z+PU0BDP3ivhe7BPSYsIldtnRrfnuMs3didUDOSa8pwPW6ATnZpew31BI
4QKUvdbDgachMwhf0qxtqC/Qd66lpMZaPmYdBFsmX5knNQ2BF1VySIYmvlfTe3l1
LnMVmLkSOX9RAVjJmbHSG4pOBWN5/FqV8k+lAw0UYuIbMk1Es0YfBbZGE3bPC5QO
v8ANCO1VbFr35s+91LmeSkbxPI6/SLnJkfGFqVsX/BcZ+opwZvjFuUeLFuIgB1tX
p28gTGhEYJldYFdYtDoBuZhLPWSB14nDG7h4ISetVxeciEYES2b3+gU5S763cms1
W+fa3JJK1eJOBYjgdV5OmiR7Bv1IUKQf5fFIoJjuKshEW9TLlEMbQ7XyvX8ZErH1
gTKdrmeGz04SBHPdIPjbp7UHqn65NaMZsrfxlI6Z/QMQ+ptxGBlzWa7S9lYDNYYs
SZIi3pqiFoJpXAbuhSQlXuFWQw0HFHoxnvrzt/e3walmfIMc+c6vT9Jq8QAoLABN
1R2wDzkZDFwFPvqjgxB59UOZoX3sY+mOxLDbKJWKLHxWow2Jkdlz7ictHViSaeS4
uWbSZyGNsQ1fbQNyePNjUYyhAGLOPJYI5oeD52QCjSZEawfawNgBp5oISRzM0wR4
cnSNgtENlichSoBwZykpTV4YfnJDIiYkaUFm4DSsccAPbbKeJ5MBw/1Gj0LtORe0
zabRNdZ+OZmHOAbtk20ZUp8TyoxddHd87gS0gHB0t7sDE97D67qytk0mojJfhc6f
Q1nKhkMmPkeLwKqIYmYOc+dMNiJHvgK0fmAAhOt+LKNwNS4aHvvXUr3Pe8KnwvL1
LIDXOvJF+GpuEmhB17b5awSVP152uhJryN589zU0J8OFtKAjs42RJtIe9tdgBxsp
FTYE7w3h0hftWM7Y/TrthKTB/P+hhWm0LtylA5VwdRoLwMaYV9PKbEMx62fKfccA
7bYa8Yg7SPGq/gBhjcoRICWwYgEetZbKSlI665GSKdGN0yohWn5s+eny+jj6B+re
rr0bz8Tcmq6dF9aKp2RPof+s2tVeM8EXmMRICv5EmQz07njyvU3gBYgLdQVCsyoM
YSXM1C1LmXQhVf8c1/R8fVSZGtg/9fOzfRXWaC8S6yp9rw/vU3syt959jJRS7Xmu
nNeEfMuKsZOzwwntyPsK8z7UgVHzVRlMpzann0avPxVVgVuHmsYIYU0r4RHOfKq6
Dmusqrhew4ALCgllujDmafjm6umYHG5D9ACuDQj0uWCu6kmSZFHYzLSBVHMkGWLv
6XxWdGwqW4VcPUltZKaD+ywUtkUwiN2rkY3txKLnwPsBHhV5oUC72XhNCbeA90f+
hOEULwBjpnraLipfLFGt4J7dHn3+thCAqx+Lm75G+NIzmQmovR+eaUFbuw+As3R3
glR2QC1FftWQu7zzmoVbH6b3Qa70xtHFCHQAkZJDMT74ChHncWE98sQlK1OOeDo5
/tjPSfBIq6KY3TNv2vK0omrXSzZKWUOZQmfKgtTnhVi3wzRL8kbWfWvamufgULy7
WZ0iaKnIkw7ahpIDMPoUniNSCs7OfKX5ZHAXGOuk7x8dubdHD2KUJrPuFKDerMbD
GKL/XSvcaX/0TmbPchzV5vVodYbMms2WyP5LlGxNC8X7+q1mWXQYlGIDq/sYWDS8
yTQ/swzaeVSndOjaJZ339qg37kT8laaB8sFgAKBwVT8+OBBxxSinwBZENqpEOhn8
CZANo9mep/hTKDA57DqI0Z5BmXerBd6DVzBmcpOOoWzmaFcB43ncyNgQwE2LQ1cO
UskrBHZjaIMbSxFHdGp8ifguGlGLbX4r5pDMuhKcZZSJLi5XvtXAr/pGBp18piEw
3daj0PJ2T8PsWCOp5gt3lUIUrgkDvIOKKJkbdbOij5O2Ucy9hqf2CTF0Xv/0NSpg
KYZEBQC9usRn/y4RR6Vos7g8TwjWLpCUddsGixyfae4yEFREhi3ABhRIdjO8JIed
8EyNWSJm/ch4A5Rv38pqCdU00f4wluq/48BLf4Wca+OXiUzz5NFfqAsdrG2fvI0t
yhOrLK6yUopBcNHus38SC3dG1pfFxhKYB3uPiNSQJO5exD6RiMbOiQiaPbaCbsST
i16W3zn7QGa2euFxP2/tHKqmTt7OddMzxXxy0M1GlYUU1nMtVkaO3gw3aev7qGV9
ckdd0nky28/ByMC/xQKERdEXdVGz04/+EXY1xhLYWuWw273Yf4dKYrFLx5ffDqb7
NYep1+YDtLNeYFauhDKNCL/awcwebLb3lAGOcDb9H3eB+OnIT+fGdTc8LGveqTZq
PRIlP0+S51MFjLpuiMp7j0JO8iMiuzMizV6MzwepEjgHHGTdXbRrpdsw7zZT0AW3
v5vfN85f1culvQIEN5CLsgHfYn5XrQkNw6sibzRmSX6rSne++6Ttxu91oJwdCwzT
GQbaaduoQc7uq9T83Ab9WJEpuIVIHi4+vTPoMznRtIAxZr8S4jRqOd1/OyExM8N5
zaMtYAFzJl0iJHsbzFSG3hJnqh+91Kq2T7DttDfqsYsurXgSTYTzvOlyWLeXJjeb
lyDvVzVS+/A0F4G81YGNJELvzhZ6YFqAjF2Ppjjr4esWF4OWl7vRmIaXjXmte1um
gNn3trw2BDIPf6TMHnZ1SXmmC+wUNI+GfMUFRnuxNGs5CO8mLiwdgH4xELS4SjjY
BAXqVg8xnJgQIBVTz34TFcU+HvuAP0BLORQPlcaUlerCxjoYBpMZcoXVUi2lk3au
W4WApPwABX494mGEt+DuNPbprnzyKy1HJwsIIrxWUsogIt+N/LmLj+PMnX2yW0SW
hUdX2k5fa1sNoSttLanRgBpJn+ZCiTfHQVWheE9gE4u8CT2Ok3K0KVgHBb2EvAmk
Gs3WsaPtKxOcQQa/Gm26+TJpqWIDNcfEkpd2rmeqVaPnl8l5BvUspo7EMcFe3mKQ
mtTp7CrG+q/HRVohnqvzowi+1THitw/ouoLKn/miTtI/SfEj88/mNc+qF06iL5+v
Qu/RSblgZf0aZuumdEIaYJNwuSNu8DO+NQblM/NGhWHtPUKBjBhruJ+5SXX36OZF
XRS2wG0kmqUESj+EPNp/9eexIkEHyMqdbNbVCuyASVqXd/YCNuz3qIN+68Y+Nela
XSaApUJQ9aIFgxrBHWPNst2dqFR1BxPbU0t7G4kfxLGk0xcHt86vuy2lKohs12NI
LNqq/x8fBeUX419F8PpjtLMZ53ei304eYgbxRrY9GVpLRuzYCzPBfL3BaOjsOiUn
V237KYbgLpqlocJlvDxFlhdclck+izM7RpmF5MiqYoi4kB8rBCOdjU7W+M33lcfT
aj+EXbcWyCr5+jji5CifssI65mEqjMB9vlplYr4RFGaSpA/pUM1QZQ3ymmGWTpwy
euvTNs6W+U4b/B3YJ12MmX17kiIsGWf9WY3Xi//dSrcI8W3zE3/NFyLH2fia4JfH
Q8KW5z0M88ZZc2KiUod0jzcOBC930MFXVL4BddTY8A8ZLnC7uhDXB4aaZFRe/AUh
TvNH+02+M622LQ26dr6zylpBBW9xcCwy0hGQSkPXpfXIGzP0kEZ1vgnDAwAFgWOe
6i3JlgyKsw4QcHvvGcBlSX5mGnM125A4nmAD4IJCDC009JWQQgzLTm71p8YMsHE3
YYaKmkJ/i9PfR21Az2KGdtbY2TAbKA0ZRBYUesc3kjYXvxVlynEelNWOODdONQck
RzLNWHV5Ym2BUwoa1mgYo2LuZSfe0OElfT8NdtxmixhzA3LvngVDqymQJhs6zYGN
61EHn2y1G8g7m7JUGxOeAtjUFlWoKfhxqzftJYgAbiOdCqJCKaYjFzCY0oOj037k
rR8V4A6BnnVe7la45e71O0FnCfUo/esfK4kME9vJs02gcUwG4rsgFvzb2PVPtnyq
aBDR/N2YFF4yNPLCsp/82ygfK9LBBHl2+l867Oh/cjpdUqJ5DiYIp/9Ao7XJms8z
DiCJm7skvhnM+UpNYYeFuoVcje2FrkJQzbrPv1doCeKyr7fPEZk1biTZDWb+6XI+
0/JENKfMGWXHW3Ey8dw8zAqpzt5lb34dRp5s0UjtYGUM5D+vVZXXukSyYpIJ++4R
ywYuwXouI6ERMw735a150YeVPPwEe6E9sDEHnLcOcptZgqopIQANF4AmE7sS79GY
fVOE+dG+9LMDGJq+myrkR1wgfDZZCYjDhqdZFbVT6zy7jmEX1Dnch0PLKzK8UAhF
jKc0bqL7V9SAtIwFN4GCqe1INxrFXoMGiE0nLQDuDjkAedU8sWszR5IlA4WOIcdP
8n5vfnr1u+4bSyDPHIHbOLnmFy1EhNYamPEzY2lqLgWHkcnh/ZE/M/aV0tmSjj9y
SszK9k1BnCUnFJ5Ge9PAO3/fk2VPe5AhsxhteTInbPNnsm24EkOGnUT76PXxXcg6
VzOqEF5X6Whx8fxV+xXAHKezUWcK9kq3z4RUomHXHxvXeUFOiqkLu8TF6OCMIUyT
CEpjWUhtq/7e99hngJx1csl+MNFqN+azvO8sSc+D2nlGcReUxpccuCXloBv2BO0h
l4C2G2XpEIvVV9QZankwXwyNdZj1qMYcKmt/khokotgxp9t7J4eKw1fMnSHzkECZ
ANcYgC2RIM08I32Q7N/L8251CH9dyKeusDArjHqcy9FmHr1+hotHvfmAXh5JX02w
4AOmtqy4NSG4SiBmZlbxuPbFm4zHw9HrV9+9oTN3h4Ov3tDFVAXjaJmRCM2l3Ti9
bE/XgAKoDaTvg2TrrlVo49X9fhnNpl4feLQGXfRzkj+VpBCOk461ipvdjARdCeWA
pMksr5ENB8bj2pKEvaVjRnhg7KPAX460ae27NiyVAasvE7RopTdf8kUaTI2/nMFR
MpVAfA5r0UU5RrMaRgQwzGEHffAGL3QCYZjFSEGlDtb5WmSsM7JP4VCNUL74YL/m
E/1IP2SO79tB1AIy3jUSVpNF7WOcCsQXxkX7s9qVINRQB46lDa7ncglnINjmSF/0
N6nt1TQdAChvPwHl1kJyF5P48KeAX2yJiFwgbBOlOEP8ne+1gh+TK9ZeM2EpJ+Ly
HIHTzYyItO1oxrp+Ie5pxQOU21UutAHr6Ce7F1BDrwuYXLU07IPHk0KDsAIkeEGa
sA5/iYj4fwqq2PWNTylKzJakSip84cBWr9g4LbDvko/RGm1H91OzohTBoa7/4u7U
Em5mXAapC43bHqzqKUeWw1dJWpcj+IN/E6JDFJjD/T7cfxjYW32r7dbdnYK8wN53
dhk3wlW/kjEC1AmTuAEwnD7a4TNAnLXc0za/eGwLQ5VJTfKI1DRPX3Gn6kJTwSB5
eO5WsLX4efqYrM1FSfv57VHy2dln+UEICowBxyMxwvR9Zjj4F3gUe3EAknIskl5T
EyQB9Ko3FlLdJ2I04Chvk2cGoIJOL5SV5IP4BHo+ucX1j4IzTTWj+CHt5XBwsHN9
LymjMubOAhOGSAto7T3TCf3dyozJJ+kKeMDhlHwVme8y3qhb63Adn5p0rdX3GU1E
H87FCszO+aNAMMKT6xT+icerfh5y1YLWIwnDgXPqoD8yJ7urfxpykPFDfQ+t2KV2
udnSfiWP/yiIR+UpgBC6PHn3HmQ8edOF75HLHwF1cdfi/KgfjDjLeyq0+aPeG1Z+
CJDoLl0G1fFBc0nSduPAwFdmjODBnESrlroB30U7ClGix+p2/o/HufPHXRc6ZRLe
UtLstdtccl38BdTU4FKvwGq7emV/wV9KjWUcpuaPx2s/acA3lidNRG05QDgiC60f
1ySYksU70Y49s5sxIqOvr3H5Tr0pg836d0QewRI65JP0Y+8+gye6KmMQYZv92diA
I692ymVGWWI5pXiy0xsWaMaiK6VLaKFmQbCifoz6C4rfGS2dai8+1mipRhTfm7xW
0pTmzIMvP6wgFF9XeYdMJIWac8w2FrilXi+4B+oY9zlusiweYyFCYdPKaWm1yFjh
LZvv9R6UITNYrGedhH73SJ1RTZ5n/pD42UvxogqOJjt1zhBEn9R34kDQgem0tcC+
vvruxS5FA/Dm3Ue/w8EDQbSYjBr92ZB7VaCWJ1p0E8V62HudH3E4kV55wvGrR6o6
AInfn2DQheqkUsu81tttyxNEfIUz0RMA6gEN012N6+HrFoznFo4ZOZkoYky6xjS0
jTF7W3pwCDReLdlHWjUlcTmmsg9oadetJddzyFQXfPyi4Endx00zyJXDGy8JNqaH
UUn5LiGzdEwtvYLu5jjbwrwpMEPAJZNJ6rkqn3b2YBtZXYcGFUoSiBzhBG84kNK7
WLHZIbCB0uwOErFc9xq450314a8FEmbgoljEMJfHYDSPfC8ZHpoPghBNyG7DUfQx
Sqx1Ke9aXzOMTn459xbohDIE6nwo9wUbzAzejIPJ34Qnf6b0YbmZLuZFJxbBwTIs
E8PWczGhPRaaJcWgUDtmOQTldOBsg33PGJtikkHFhxCUMY4AztlLLoke+Wpv/3uE
`pragma protect end_protected
