-- MebX_Qsys_Project_Burst_tb.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity MebX_Qsys_Project_Burst_tb is
end entity MebX_Qsys_Project_Burst_tb;

architecture rtl of MebX_Qsys_Project_Burst_tb is
	component MebX_Qsys_Project_Burst is
		port (
			clk100_clk                       : in  std_logic := 'X'; -- clk
			clk200_clk                       : in  std_logic := 'X'; -- clk
			clk50_clk                        : in  std_logic := 'X'; -- clk
			comm_a_conduit_end_spw_si_signal : in  std_logic := 'X'; -- spw_si_signal
			comm_a_conduit_end_spw_di_signal : in  std_logic := 'X'; -- spw_di_signal
			comm_a_conduit_end_spw_do_signal : out std_logic;        -- spw_do_signal
			comm_a_conduit_end_spw_so_signal : out std_logic;        -- spw_so_signal
			rst_reset_n                      : in  std_logic := 'X'; -- reset_n
			timer_1ms_external_port_export   : out std_logic;        -- export
			timer_1us_external_port_export   : out std_logic         -- export
		);
	end component MebX_Qsys_Project_Burst;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_conduit_bfm is
		port (
			clk               : in  std_logic                    := 'X';             -- clk
			sig_spw_si_signal : out std_logic_vector(0 downto 0);                    -- spw_si_signal
			sig_spw_di_signal : out std_logic_vector(0 downto 0);                    -- spw_di_signal
			sig_spw_do_signal : in  std_logic_vector(0 downto 0) := (others => 'X'); -- spw_do_signal
			sig_spw_so_signal : in  std_logic_vector(0 downto 0) := (others => 'X'); -- spw_so_signal
			reset             : in  std_logic                    := 'X'              -- reset
		);
	end component altera_conduit_bfm;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_conduit_bfm_0002 is
		port (
			sig_export : in std_logic_vector(0 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0002;

	signal mebx_qsys_project_burst_inst_clk100_bfm_clk_clk                           : std_logic;                    -- MebX_Qsys_Project_Burst_inst_clk100_bfm:clk -> [MebX_Qsys_Project_Burst_inst:clk100_clk, MebX_Qsys_Project_Burst_inst_comm_a_conduit_end_bfm:clk, MebX_Qsys_Project_Burst_inst_rst_bfm:clk]
	signal mebx_qsys_project_burst_inst_clk200_bfm_clk_clk                           : std_logic;                    -- MebX_Qsys_Project_Burst_inst_clk200_bfm:clk -> MebX_Qsys_Project_Burst_inst:clk200_clk
	signal mebx_qsys_project_burst_inst_clk50_bfm_clk_clk                            : std_logic;                    -- MebX_Qsys_Project_Burst_inst_clk50_bfm:clk -> MebX_Qsys_Project_Burst_inst:clk50_clk
	signal mebx_qsys_project_burst_inst_comm_a_conduit_end_spw_do_signal             : std_logic;                    -- MebX_Qsys_Project_Burst_inst:comm_a_conduit_end_spw_do_signal -> MebX_Qsys_Project_Burst_inst_comm_a_conduit_end_bfm:sig_spw_do_signal
	signal mebx_qsys_project_burst_inst_comm_a_conduit_end_spw_so_signal             : std_logic;                    -- MebX_Qsys_Project_Burst_inst:comm_a_conduit_end_spw_so_signal -> MebX_Qsys_Project_Burst_inst_comm_a_conduit_end_bfm:sig_spw_so_signal
	signal mebx_qsys_project_burst_inst_comm_a_conduit_end_bfm_conduit_spw_di_signal : std_logic_vector(0 downto 0); -- MebX_Qsys_Project_Burst_inst_comm_a_conduit_end_bfm:sig_spw_di_signal -> MebX_Qsys_Project_Burst_inst:comm_a_conduit_end_spw_di_signal
	signal mebx_qsys_project_burst_inst_comm_a_conduit_end_bfm_conduit_spw_si_signal : std_logic_vector(0 downto 0); -- MebX_Qsys_Project_Burst_inst_comm_a_conduit_end_bfm:sig_spw_si_signal -> MebX_Qsys_Project_Burst_inst:comm_a_conduit_end_spw_si_signal
	signal mebx_qsys_project_burst_inst_timer_1ms_external_port_export               : std_logic;                    -- MebX_Qsys_Project_Burst_inst:timer_1ms_external_port_export -> MebX_Qsys_Project_Burst_inst_timer_1ms_external_port_bfm:sig_export
	signal mebx_qsys_project_burst_inst_timer_1us_external_port_export               : std_logic;                    -- MebX_Qsys_Project_Burst_inst:timer_1us_external_port_export -> MebX_Qsys_Project_Burst_inst_timer_1us_external_port_bfm:sig_export
	signal mebx_qsys_project_burst_inst_rst_bfm_reset_reset                          : std_logic;                    -- MebX_Qsys_Project_Burst_inst_rst_bfm:reset -> MebX_Qsys_Project_Burst_inst:rst_reset_n

begin

	mebx_qsys_project_burst_inst : component MebX_Qsys_Project_Burst
		port map (
			clk100_clk                       => mebx_qsys_project_burst_inst_clk100_bfm_clk_clk,                              --                  clk100.clk
			clk200_clk                       => mebx_qsys_project_burst_inst_clk200_bfm_clk_clk,                              --                  clk200.clk
			clk50_clk                        => mebx_qsys_project_burst_inst_clk50_bfm_clk_clk,                               --                   clk50.clk
			comm_a_conduit_end_spw_si_signal => mebx_qsys_project_burst_inst_comm_a_conduit_end_bfm_conduit_spw_si_signal(0), --      comm_a_conduit_end.spw_si_signal
			comm_a_conduit_end_spw_di_signal => mebx_qsys_project_burst_inst_comm_a_conduit_end_bfm_conduit_spw_di_signal(0), --                        .spw_di_signal
			comm_a_conduit_end_spw_do_signal => mebx_qsys_project_burst_inst_comm_a_conduit_end_spw_do_signal,                --                        .spw_do_signal
			comm_a_conduit_end_spw_so_signal => mebx_qsys_project_burst_inst_comm_a_conduit_end_spw_so_signal,                --                        .spw_so_signal
			rst_reset_n                      => mebx_qsys_project_burst_inst_rst_bfm_reset_reset,                             --                     rst.reset_n
			timer_1ms_external_port_export   => mebx_qsys_project_burst_inst_timer_1ms_external_port_export,                  -- timer_1ms_external_port.export
			timer_1us_external_port_export   => mebx_qsys_project_burst_inst_timer_1us_external_port_export                   -- timer_1us_external_port.export
		);

	mebx_qsys_project_burst_inst_clk100_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 100000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => mebx_qsys_project_burst_inst_clk100_bfm_clk_clk  -- clk.clk
		);

	mebx_qsys_project_burst_inst_clk200_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 200000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => mebx_qsys_project_burst_inst_clk200_bfm_clk_clk  -- clk.clk
		);

	mebx_qsys_project_burst_inst_clk50_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => mebx_qsys_project_burst_inst_clk50_bfm_clk_clk  -- clk.clk
		);

	mebx_qsys_project_burst_inst_comm_a_conduit_end_bfm : component altera_conduit_bfm
		port map (
			clk                  => mebx_qsys_project_burst_inst_clk100_bfm_clk_clk,                           --     clk.clk
			sig_spw_si_signal    => mebx_qsys_project_burst_inst_comm_a_conduit_end_bfm_conduit_spw_si_signal, -- conduit.spw_si_signal
			sig_spw_di_signal    => mebx_qsys_project_burst_inst_comm_a_conduit_end_bfm_conduit_spw_di_signal, --        .spw_di_signal
			sig_spw_do_signal(0) => mebx_qsys_project_burst_inst_comm_a_conduit_end_spw_do_signal,             --        .spw_do_signal
			sig_spw_so_signal(0) => mebx_qsys_project_burst_inst_comm_a_conduit_end_spw_so_signal,             --        .spw_so_signal
			reset                => '0'                                                                        -- (terminated)
		);

	mebx_qsys_project_burst_inst_rst_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => mebx_qsys_project_burst_inst_rst_bfm_reset_reset, -- reset.reset_n
			clk   => mebx_qsys_project_burst_inst_clk100_bfm_clk_clk   --   clk.clk
		);

	mebx_qsys_project_burst_inst_timer_1ms_external_port_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export(0) => mebx_qsys_project_burst_inst_timer_1ms_external_port_export  -- conduit.export
		);

	mebx_qsys_project_burst_inst_timer_1us_external_port_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export(0) => mebx_qsys_project_burst_inst_timer_1us_external_port_export  -- conduit.export
		);

end architecture rtl; -- of MebX_Qsys_Project_Burst_tb
