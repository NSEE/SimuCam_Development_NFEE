library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity windowing_machine_ent is
	port(
		clk_i : in std_logic;
		rst_i : in std_logic
	);
end entity windowing_machine_ent;

architecture RTL of windowing_machine_ent is
	
begin

end architecture RTL;
