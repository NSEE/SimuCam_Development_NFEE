// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.



// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// $Id: //acds/rel/18.1std/ip/merlin/altera_merlin_router/altera_merlin_router.sv.terp#1 $
// $Revision: #1 $
// $Date: 2018/07/18 $
// $Author: psgswbuild $

// -------------------------------------------------------
// Merlin Router
//
// Asserts the appropriate one-hot encoded channel based on 
// either (a) the address or (b) the dest id. The DECODER_TYPE
// parameter controls this behaviour. 0 means address decoder,
// 1 means dest id decoder.
//
// In the case of (a), it also sets the destination id.
// -------------------------------------------------------

`timescale 1 ns / 1 ns

module MebX_Qsys_Project_mm_interconnect_0_router_004_default_decode
  #(
     parameter DEFAULT_CHANNEL = 1,
               DEFAULT_WR_CHANNEL = -1,
               DEFAULT_RD_CHANNEL = -1,
               DEFAULT_DESTID = 29 
   )
  (output [367 - 362 : 0] default_destination_id,
   output [34-1 : 0] default_wr_channel,
   output [34-1 : 0] default_rd_channel,
   output [34-1 : 0] default_src_channel
  );

  assign default_destination_id = 
    DEFAULT_DESTID[367 - 362 : 0];

  generate
    if (DEFAULT_CHANNEL == -1) begin : no_default_channel_assignment
      assign default_src_channel = '0;
    end
    else begin : default_channel_assignment
      assign default_src_channel = 34'b1 << DEFAULT_CHANNEL;
    end
  endgenerate

  generate
    if (DEFAULT_RD_CHANNEL == -1) begin : no_default_rw_channel_assignment
      assign default_wr_channel = '0;
      assign default_rd_channel = '0;
    end
    else begin : default_rw_channel_assignment
      assign default_wr_channel = 34'b1 << DEFAULT_WR_CHANNEL;
      assign default_rd_channel = 34'b1 << DEFAULT_RD_CHANNEL;
    end
  endgenerate

endmodule


module MebX_Qsys_Project_mm_interconnect_0_router_004
(
    // -------------------
    // Clock & Reset
    // -------------------
    input clk,
    input reset,

    // -------------------
    // Command Sink (Input)
    // -------------------
    input                       sink_valid,
    input  [381-1 : 0]    sink_data,
    input                       sink_startofpacket,
    input                       sink_endofpacket,
    output                      sink_ready,

    // -------------------
    // Command Source (Output)
    // -------------------
    output                          src_valid,
    output reg [381-1    : 0] src_data,
    output reg [34-1 : 0] src_channel,
    output                          src_startofpacket,
    output                          src_endofpacket,
    input                           src_ready
);

    // -------------------------------------------------------
    // Local parameters and variables
    // -------------------------------------------------------
    localparam PKT_ADDR_H = 321;
    localparam PKT_ADDR_L = 288;
    localparam PKT_DEST_ID_H = 367;
    localparam PKT_DEST_ID_L = 362;
    localparam PKT_PROTECTION_H = 371;
    localparam PKT_PROTECTION_L = 369;
    localparam ST_DATA_W = 381;
    localparam ST_CHANNEL_W = 34;
    localparam DECODER_TYPE = 0;

    localparam PKT_TRANS_WRITE = 324;
    localparam PKT_TRANS_READ  = 325;

    localparam PKT_ADDR_W = PKT_ADDR_H-PKT_ADDR_L + 1;
    localparam PKT_DEST_ID_W = PKT_DEST_ID_H-PKT_DEST_ID_L + 1;



    // -------------------------------------------------------
    // Figure out the number of bits to mask off for each slave span
    // during address decoding
    // -------------------------------------------------------
    localparam PAD0 = log2ceil(64'h80000000 - 64'h0); 
    localparam PAD1 = log2ceil(64'h100002000 - 64'h100000000); 
    localparam PAD2 = log2ceil(64'h10000a000 - 64'h100008000); 
    localparam PAD3 = log2ceil(64'h100012000 - 64'h100010000); 
    localparam PAD4 = log2ceil(64'h10001a000 - 64'h100018000); 
    localparam PAD5 = log2ceil(64'h100022000 - 64'h100020000); 
    localparam PAD6 = log2ceil(64'h10002a000 - 64'h100028000); 
    localparam PAD7 = log2ceil(64'h100032000 - 64'h100030000); 
    localparam PAD8 = log2ceil(64'h10003a000 - 64'h100038000); 
    localparam PAD9 = log2ceil(64'h100042000 - 64'h100040000); 
    localparam PAD10 = log2ceil(64'h10004a000 - 64'h100048000); 
    localparam PAD11 = log2ceil(64'h100052000 - 64'h100050000); 
    localparam PAD12 = log2ceil(64'h10005a000 - 64'h100058000); 
    localparam PAD13 = log2ceil(64'h200008000 - 64'h200000000); 
    // -------------------------------------------------------
    // Work out which address bits are significant based on the
    // address range of the slaves. If the required width is too
    // large or too small, we use the address field width instead.
    // -------------------------------------------------------
    localparam ADDR_RANGE = 64'h200008000;
    localparam RANGE_ADDR_WIDTH = log2ceil(ADDR_RANGE);
    localparam OPTIMIZED_ADDR_H = (RANGE_ADDR_WIDTH > PKT_ADDR_W) ||
                                  (RANGE_ADDR_WIDTH == 0) ?
                                        PKT_ADDR_H :
                                        PKT_ADDR_L + RANGE_ADDR_WIDTH - 1;

    localparam RG = RANGE_ADDR_WIDTH-1;
    localparam REAL_ADDRESS_RANGE = OPTIMIZED_ADDR_H - PKT_ADDR_L;

      reg [PKT_ADDR_W-1 : 0] address;
      always @* begin
        address = {PKT_ADDR_W{1'b0}};
        address [REAL_ADDRESS_RANGE:0] = sink_data[OPTIMIZED_ADDR_H : PKT_ADDR_L];
      end   

    // -------------------------------------------------------
    // Pass almost everything through, untouched
    // -------------------------------------------------------
    assign sink_ready        = src_ready;
    assign src_valid         = sink_valid;
    assign src_startofpacket = sink_startofpacket;
    assign src_endofpacket   = sink_endofpacket;
    wire [PKT_DEST_ID_W-1:0] default_destid;
    wire [34-1 : 0] default_src_channel;




    // -------------------------------------------------------
    // Write and read transaction signals
    // -------------------------------------------------------
    wire write_transaction;
    assign write_transaction = sink_data[PKT_TRANS_WRITE];


    MebX_Qsys_Project_mm_interconnect_0_router_004_default_decode the_default_decode(
      .default_destination_id (default_destid),
      .default_wr_channel   (),
      .default_rd_channel   (),
      .default_src_channel  (default_src_channel)
    );

    always @* begin
        src_data    = sink_data;
        src_channel = default_src_channel;
        src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = default_destid;

        // --------------------------------------------------
        // Address Decoder
        // Sets the channel and destination ID based on the address
        // --------------------------------------------------

    // ( 0x0 .. 0x80000000 )
    if ( {address[RG:PAD0],{PAD0{1'b0}}} == 34'h0   ) begin
            src_channel = 34'b00000000000010;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 29;
    end

    // ( 0x100000000 .. 0x100002000 )
    if ( {address[RG:PAD1],{PAD1{1'b0}}} == 34'h100000000  && write_transaction  ) begin
            src_channel = 34'b00000000000100;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 0;
    end

    // ( 0x100008000 .. 0x10000a000 )
    if ( {address[RG:PAD2],{PAD2{1'b0}}} == 34'h100008000  && write_transaction  ) begin
            src_channel = 34'b00000100000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 1;
    end

    // ( 0x100010000 .. 0x100012000 )
    if ( {address[RG:PAD3],{PAD3{1'b0}}} == 34'h100010000  && write_transaction  ) begin
            src_channel = 34'b00000000001000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 3;
    end

    // ( 0x100018000 .. 0x10001a000 )
    if ( {address[RG:PAD4],{PAD4{1'b0}}} == 34'h100018000  && write_transaction  ) begin
            src_channel = 34'b00001000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 4;
    end

    // ( 0x100020000 .. 0x100022000 )
    if ( {address[RG:PAD5],{PAD5{1'b0}}} == 34'h100020000  && write_transaction  ) begin
            src_channel = 34'b00000000010000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 6;
    end

    // ( 0x100028000 .. 0x10002a000 )
    if ( {address[RG:PAD6],{PAD6{1'b0}}} == 34'h100028000  && write_transaction  ) begin
            src_channel = 34'b00010000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 7;
    end

    // ( 0x100030000 .. 0x100032000 )
    if ( {address[RG:PAD7],{PAD7{1'b0}}} == 34'h100030000  && write_transaction  ) begin
            src_channel = 34'b00000000100000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 9;
    end

    // ( 0x100038000 .. 0x10003a000 )
    if ( {address[RG:PAD8],{PAD8{1'b0}}} == 34'h100038000  && write_transaction  ) begin
            src_channel = 34'b00100000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 10;
    end

    // ( 0x100040000 .. 0x100042000 )
    if ( {address[RG:PAD9],{PAD9{1'b0}}} == 34'h100040000  && write_transaction  ) begin
            src_channel = 34'b00000001000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 12;
    end

    // ( 0x100048000 .. 0x10004a000 )
    if ( {address[RG:PAD10],{PAD10{1'b0}}} == 34'h100048000  && write_transaction  ) begin
            src_channel = 34'b01000000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 13;
    end

    // ( 0x100050000 .. 0x100052000 )
    if ( {address[RG:PAD11],{PAD11{1'b0}}} == 34'h100050000  && write_transaction  ) begin
            src_channel = 34'b00000010000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 15;
    end

    // ( 0x100058000 .. 0x10005a000 )
    if ( {address[RG:PAD12],{PAD12{1'b0}}} == 34'h100058000  && write_transaction  ) begin
            src_channel = 34'b10000000000000;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 16;
    end

    // ( 0x200000000 .. 0x200008000 )
    if ( {address[RG:PAD13],{PAD13{1'b0}}} == 34'h200000000   ) begin
            src_channel = 34'b00000000000001;
            src_data[PKT_DEST_ID_H:PKT_DEST_ID_L] = 19;
    end

end


    // --------------------------------------------------
    // Ceil(log2()) function
    // --------------------------------------------------
    function integer log2ceil;
        input reg[65:0] val;
        reg [65:0] i;

        begin
            i = 1;
            log2ceil = 0;

            while (i < val) begin
                log2ceil = log2ceil + 1;
                i = i << 1;
            end
        end
    endfunction

endmodule


