library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity avalon_buffer_R_stimuli is
	generic(
		g_ADDRESS_WIDTH : natural range 1 to 64;
		g_DATA_WIDTH    : natural range 1 to 256
	);
	port(
		clk_i                   : in  std_logic;
		rst_i                   : in  std_logic;
		avalon_mm_waitrequest_i : in  std_logic; --                                     -- avalon_mm.waitrequest
		avalon_mm_address_o     : out std_logic_vector((g_ADDRESS_WIDTH - 1) downto 0); --          .address
		avalon_mm_write_o       : out std_logic; --                                     --          .write
		avalon_mm_writedata_o   : out std_logic_vector((g_DATA_WIDTH - 1) downto 0) --  --          .writedata
	);
end entity avalon_buffer_R_stimuli;

architecture RTL of avalon_buffer_R_stimuli is
	-- ccd image data
	constant c_CCD_IMGDATA_LENGTH : natural                                       := 4352;
	signal s_ccd_imgdata_cnt      : natural range 0 to (c_CCD_IMGDATA_LENGTH - 1) := 0;
	type t_ccd_imgdata is array (0 to (c_CCD_IMGDATA_LENGTH - 1)) of std_logic_vector(255 downto 0);
	constant c_CCD_IMGDATA        : t_ccd_imgdata                                 := (
		x"000F000E000D000C000B000A0009000800070006000500040003000200010000",
		x"001F001E001D001C001B001A0019001800170016001500140013001200110010",
		x"002F002E002D002C002B002A0029002800270026002500240023002200210020",
		x"003F003E003D003C003B003A0039003800370036003500340033003200310030",
		x"004B004A0049004800470046004500440043004200410040FFFFFFFFFFFFFFFE",
		x"005B005A0059005800570056005500540053005200510050004F004E004D004C",
		x"006B006A0069006800670066006500640063006200610060005F005E005D005C",
		x"007B007A0079007800770076007500740073007200710070006F006E006D006C",
		x"00870086008500840083008200810080FFFFFFFFFFFFFFFF007F007E007D007C",
		x"00970096009500940093009200910090008F008E008D008C008B008A00890088",
		x"00A700A600A500A400A300A200A100A0009F009E009D009C009B009A00990098",
		x"00B700B600B500B400B300B200B100B000AF00AE00AD00AC00AB00AA00A900A8",
		x"00C300C200C100C0FFFFFFFFFFFFFFFF00BF00BE00BD00BC00BB00BA00B900B8",
		x"00D300D200D100D000CF00CE00CD00CC00CB00CA00C900C800C700C600C500C4",
		x"00E300E200E100E000DF00DE00DD00DC00DB00DA00D900D800D700D600D500D4",
		x"00F300F200F100F000EF00EE00ED00EC00EB00EA00E900E800E700E600E500E4",
		x"FFFFFFFFFFFFFFFF00FF00FE00FD00FC00FB00FA00F900F800F700F600F500F4",
		x"010F010E010D010C010B010A0109010801070106010501040103010201010100",
		x"011F011E011D011C011B011A0119011801170116011501140113011201110110",
		x"012F012E012D012C012B012A0129012801270126012501240123012201210120",
		x"013F013E013D013C013B013A0139013801370136013501340133013201310130",
		x"014B014A0149014801470146014501440143014201410140FFFFFFFFFFFFFFFF",
		x"015B015A0159015801570156015501540153015201510150014F014E014D014C",
		x"016B016A0169016801670166016501640163016201610160015F015E015D015C",
		x"017B017A0179017801770176017501740173017201710170016F016E016D016C",
		x"01870186018501840183018201810180FFFFFFFFFFFFFFFF017F017E017D017C",
		x"01970196019501940193019201910190018F018E018D018C018B018A01890188",
		x"01A701A601A501A401A301A201A101A0019F019E019D019C019B019A01990198",
		x"01B701B601B501B401B301B201B101B001AF01AE01AD01AC01AB01AA01A901A8",
		x"01C301C201C101C0FFFFFFFFFFFFFFFF01BF01BE01BD01BC01BB01BA01B901B8",
		x"01D301D201D101D001CF01CE01CD01CC01CB01CA01C901C801C701C601C501C4",
		x"01E301E201E101E001DF01DE01DD01DC01DB01DA01D901D801D701D601D501D4",
		x"01F301F201F101F001EF01EE01ED01EC01EB01EA01E901E801E701E601E501E4",
		x"FFFFFFFFFFFFFFFF01FF01FE01FD01FC01FB01FA01F901F801F701F601F501F4",
		x"020F020E020D020C020B020A0209020802070206020502040203020202010200",
		x"021F021E021D021C021B021A0219021802170216021502140213021202110210",
		x"022F022E022D022C022B022A0229022802270226022502240223022202210220",
		x"023F023E023D023C023B023A0239023802370236023502340233023202310230",
		x"024B024A0249024802470246024502440243024202410240FFFFFFFFFFFFFFFF",
		x"025B025A0259025802570256025502540253025202510250024F024E024D024C",
		x"026B026A0269026802670266026502640263026202610260025F025E025D025C",
		x"027B027A0279027802770276027502740273027202710270026F026E026D026C",
		x"02870286028502840283028202810280FFFFFFFFFFFFFFFF027F027E027D027C",
		x"02970296029502940293029202910290028F028E028D028C028B028A02890288",
		x"02A702A602A502A402A302A202A102A0029F029E029D029C029B029A02990298",
		x"02B702B602B502B402B302B202B102B002AF02AE02AD02AC02AB02AA02A902A8",
		x"02C302C202C102C0FFFFFFFFFFFFFFFF02BF02BE02BD02BC02BB02BA02B902B8",
		x"02D302D202D102D002CF02CE02CD02CC02CB02CA02C902C802C702C602C502C4",
		x"02E302E202E102E002DF02DE02DD02DC02DB02DA02D902D802D702D602D502D4",
		x"02F302F202F102F002EF02EE02ED02EC02EB02EA02E902E802E702E602E502E4",
		x"FFFFFFFFFFFFFFFF02FF02FE02FD02FC02FB02FA02F902F802F702F602F502F4",
		x"030F030E030D030C030B030A0309030803070306030503040303030203010300",
		x"031F031E031D031C031B031A0319031803170316031503140313031203110310",
		x"032F032E032D032C032B032A0329032803270326032503240323032203210320",
		x"033F033E033D033C033B033A0339033803370336033503340333033203310330",
		x"034B034A0349034803470346034503440343034203410340FFFFFFFFFFFFFFFF",
		x"035B035A0359035803570356035503540353035203510350034F034E034D034C",
		x"036B036A0369036803670366036503640363036203610360035F035E035D035C",
		x"037B037A0379037803770376037503740373037203710370036F036E036D036C",
		x"03870386038503840383038203810380FFFFFFFFFFFFFFFF037F037E037D037C",
		x"03970396039503940393039203910390038F038E038D038C038B038A03890388",
		x"03A703A603A503A403A303A203A103A0039F039E039D039C039B039A03990398",
		x"03B703B603B503B403B303B203B103B003AF03AE03AD03AC03AB03AA03A903A8",
		x"03C303C203C103C0FFFFFFFFFFFFFFFF03BF03BE03BD03BC03BB03BA03B903B8",
		x"03D303D203D103D003CF03CE03CD03CC03CB03CA03C903C803C703C603C503C4",
		x"03E303E203E103E003DF03DE03DD03DC03DB03DA03D903D803D703D603D503D4",
		x"03F303F203F103F003EF03EE03ED03EC03EB03EA03E903E803E703E603E503E4",
		x"FFFFFFFFFFFFFFFF03FF03FE03FD03FC03FB03FA03F903F803F703F603F503F4",
		x"040F040E040D040C040B040A0409040804070406040504040403040204010400",
		x"041F041E041D041C041B041A0419041804170416041504140413041204110410",
		x"042F042E042D042C042B042A0429042804270426042504240423042204210420",
		x"043F043E043D043C043B043A0439043804370436043504340433043204310430",
		x"044B044A0449044804470446044504440443044204410440FFFFFFFFFFFFFFFF",
		x"045B045A0459045804570456045504540453045204510450044F044E044D044C",
		x"046B046A0469046804670466046504640463046204610460045F045E045D045C",
		x"047B047A0479047804770476047504740473047204710470046F046E046D046C",
		x"04870486048504840483048204810480FFFFFFFFFFFFFFFF047F047E047D047C",
		x"04970496049504940493049204910490048F048E048D048C048B048A04890488",
		x"04A704A604A504A404A304A204A104A0049F049E049D049C049B049A04990498",
		x"04B704B604B504B404B304B204B104B004AF04AE04AD04AC04AB04AA04A904A8",
		x"04C304C204C104C0FFFFFFFFFFFFFFFF04BF04BE04BD04BC04BB04BA04B904B8",
		x"04D304D204D104D004CF04CE04CD04CC04CB04CA04C904C804C704C604C504C4",
		x"04E304E204E104E004DF04DE04DD04DC04DB04DA04D904D804D704D604D504D4",
		x"04F304F204F104F004EF04EE04ED04EC04EB04EA04E904E804E704E604E504E4",
		x"FFFFFFFFFFFFFFFF04FF04FE04FD04FC04FB04FA04F904F804F704F604F504F4",
		x"050F050E050D050C050B050A0509050805070506050505040503050205010500",
		x"051F051E051D051C051B051A0519051805170516051505140513051205110510",
		x"052F052E052D052C052B052A0529052805270526052505240523052205210520",
		x"053F053E053D053C053B053A0539053805370536053505340533053205310530",
		x"054B054A0549054805470546054505440543054205410540FFFFFFFFFFFFFFFF",
		x"055B055A0559055805570556055505540553055205510550054F054E054D054C",
		x"056B056A0569056805670566056505640563056205610560055F055E055D055C",
		x"057B057A0579057805770576057505740573057205710570056F056E056D056C",
		x"05870586058505840583058205810580FFFFFFFFFFFFFFFF057F057E057D057C",
		x"05970596059505940593059205910590058F058E058D058C058B058A05890588",
		x"05A705A605A505A405A305A205A105A0059F059E059D059C059B059A05990598",
		x"05B705B605B505B405B305B205B105B005AF05AE05AD05AC05AB05AA05A905A8",
		x"05C305C205C105C0FFFFFFFFFFFFFFFF05BF05BE05BD05BC05BB05BA05B905B8",
		x"05D305D205D105D005CF05CE05CD05CC05CB05CA05C905C805C705C605C505C4",
		x"05E305E205E105E005DF05DE05DD05DC05DB05DA05D905D805D705D605D505D4",
		x"05F305F205F105F005EF05EE05ED05EC05EB05EA05E905E805E705E605E505E4",
		x"FFFFFFFFFFFFFFFF05FF05FE05FD05FC05FB05FA05F905F805F705F605F505F4",
		x"060F060E060D060C060B060A0609060806070606060506040603060206010600",
		x"061F061E061D061C061B061A0619061806170616061506140613061206110610",
		x"062F062E062D062C062B062A0629062806270626062506240623062206210620",
		x"063F063E063D063C063B063A0639063806370636063506340633063206310630",
		x"064B064A0649064806470646064506440643064206410640FFFFFFFFFFFFFFFF",
		x"065B065A0659065806570656065506540653065206510650064F064E064D064C",
		x"066B066A0669066806670666066506640663066206610660065F065E065D065C",
		x"067B067A0679067806770676067506740673067206710670066F066E066D066C",
		x"06870686068506840683068206810680FFFFFFFFFFFFFFFF067F067E067D067C",
		x"06970696069506940693069206910690068F068E068D068C068B068A06890688",
		x"06A706A606A506A406A306A206A106A0069F069E069D069C069B069A06990698",
		x"06B706B606B506B406B306B206B106B006AF06AE06AD06AC06AB06AA06A906A8",
		x"06C306C206C106C0FFFFFFFFFFFFFFFF06BF06BE06BD06BC06BB06BA06B906B8",
		x"06D306D206D106D006CF06CE06CD06CC06CB06CA06C906C806C706C606C506C4",
		x"06E306E206E106E006DF06DE06DD06DC06DB06DA06D906D806D706D606D506D4",
		x"06F306F206F106F006EF06EE06ED06EC06EB06EA06E906E806E706E606E506E4",
		x"FFFFFFFFFFFFFFFF06FF06FE06FD06FC06FB06FA06F906F806F706F606F506F4",
		x"070F070E070D070C070B070A0709070807070706070507040703070207010700",
		x"071F071E071D071C071B071A0719071807170716071507140713071207110710",
		x"072F072E072D072C072B072A0729072807270726072507240723072207210720",
		x"073F073E073D073C073B073A0739073807370736073507340733073207310730",
		x"074B074A0749074807470746074507440743074207410740FFFFFFFFFFFFFFFF",
		x"075B075A0759075807570756075507540753075207510750074F074E074D074C",
		x"076B076A0769076807670766076507640763076207610760075F075E075D075C",
		x"077B077A0779077807770776077507740773077207710770076F076E076D076C",
		x"07870786078507840783078207810780FFFFFFFFFFFFFFFF077F077E077D077C",
		x"07970796079507940793079207910790078F078E078D078C078B078A07890788",
		x"07A707A607A507A407A307A207A107A0079F079E079D079C079B079A07990798",
		x"07B707B607B507B407B307B207B107B007AF07AE07AD07AC07AB07AA07A907A8",
		x"07C307C207C107C0FFFFFFFFFFFFFFFF07BF07BE07BD07BC07BB07BA07B907B8",
		x"07D307D207D107D007CF07CE07CD07CC07CB07CA07C907C807C707C607C507C4",
		x"07E307E207E107E007DF07DE07DD07DC07DB07DA07D907D807D707D607D507D4",
		x"07F307F207F107F007EF07EE07ED07EC07EB07EA07E907E807E707E607E507E4",
		x"FFFFFFFFFFFFFFFF07FF07FE07FD07FC07FB07FA07F907F807F707F607F507F4",
		x"080F080E080D080C080B080A0809080808070806080508040803080208010800",
		x"081F081E081D081C081B081A0819081808170816081508140813081208110810",
		x"082F082E082D082C082B082A0829082808270826082508240823082208210820",
		x"083F083E083D083C083B083A0839083808370836083508340833083208310830",
		x"084B084A0849084808470846084508440843084208410840FFFFFFFFFFFFFFFF",
		x"085B085A0859085808570856085508540853085208510850084F084E084D084C",
		x"086B086A0869086808670866086508640863086208610860085F085E085D085C",
		x"087B087A0879087808770876087508740873087208710870086F086E086D086C",
		x"08870886088508840883088208810880FFFFFFFFFFFFFFFF087F087E087D087C",
		x"08970896089508940893089208910890088F088E088D088C088B088A08890888",
		x"08A708A608A508A408A308A208A108A0089F089E089D089C089B089A08990898",
		x"08B708B608B508B408B308B208B108B008AF08AE08AD08AC08AB08AA08A908A8",
		x"08C308C208C108C0FFFFFFFFFFFFFFFF08BF08BE08BD08BC08BB08BA08B908B8",
		x"08D308D208D108D008CF08CE08CD08CC08CB08CA08C908C808C708C608C508C4",
		x"08E308E208E108E008DF08DE08DD08DC08DB08DA08D908D808D708D608D508D4",
		x"08F308F208F108F008EF08EE08ED08EC08EB08EA08E908E808E708E608E508E4",
		x"FFFFFFFFFFFFFFFF08FF08FE08FD08FC08FB08FA08F908F808F708F608F508F4",
		x"090F090E090D090C090B090A0909090809070906090509040903090209010900",
		x"091F091E091D091C091B091A0919091809170916091509140913091209110910",
		x"092F092E092D092C092B092A0929092809270926092509240923092209210920",
		x"093F093E093D093C093B093A0939093809370936093509340933093209310930",
		x"094B094A0949094809470946094509440943094209410940FFFFFFFFFFFFFFFF",
		x"095B095A0959095809570956095509540953095209510950094F094E094D094C",
		x"096B096A0969096809670966096509640963096209610960095F095E095D095C",
		x"097B097A0979097809770976097509740973097209710970096F096E096D096C",
		x"09870986098509840983098209810980FFFFFFFFFFFFFFFF097F097E097D097C",
		x"09970996099509940993099209910990098F098E098D098C098B098A09890988",
		x"09A709A609A509A409A309A209A109A0099F099E099D099C099B099A09990998",
		x"09B709B609B509B409B309B209B109B009AF09AE09AD09AC09AB09AA09A909A8",
		x"09C309C209C109C0FFFFFFFFFFFFFFFF09BF09BE09BD09BC09BB09BA09B909B8",
		x"09D309D209D109D009CF09CE09CD09CC09CB09CA09C909C809C709C609C509C4",
		x"09E309E209E109E009DF09DE09DD09DC09DB09DA09D909D809D709D609D509D4",
		x"09F309F209F109F009EF09EE09ED09EC09EB09EA09E909E809E709E609E509E4",
		x"FFFFFFFFFFFFFFFF09FF09FE09FD09FC09FB09FA09F909F809F709F609F509F4",
		x"0A0F0A0E0A0D0A0C0A0B0A0A0A090A080A070A060A050A040A030A020A010A00",
		x"0A1F0A1E0A1D0A1C0A1B0A1A0A190A180A170A160A150A140A130A120A110A10",
		x"0A2F0A2E0A2D0A2C0A2B0A2A0A290A280A270A260A250A240A230A220A210A20",
		x"0A3F0A3E0A3D0A3C0A3B0A3A0A390A380A370A360A350A340A330A320A310A30",
		x"0A4B0A4A0A490A480A470A460A450A440A430A420A410A40FFFFFFFFFFFFFFFF",
		x"0A5B0A5A0A590A580A570A560A550A540A530A520A510A500A4F0A4E0A4D0A4C",
		x"0A6B0A6A0A690A680A670A660A650A640A630A620A610A600A5F0A5E0A5D0A5C",
		x"0A7B0A7A0A790A780A770A760A750A740A730A720A710A700A6F0A6E0A6D0A6C",
		x"0A870A860A850A840A830A820A810A80FFFFFFFFFFFFFFFF0A7F0A7E0A7D0A7C",
		x"0A970A960A950A940A930A920A910A900A8F0A8E0A8D0A8C0A8B0A8A0A890A88",
		x"0AA70AA60AA50AA40AA30AA20AA10AA00A9F0A9E0A9D0A9C0A9B0A9A0A990A98",
		x"0AB70AB60AB50AB40AB30AB20AB10AB00AAF0AAE0AAD0AAC0AAB0AAA0AA90AA8",
		x"0AC30AC20AC10AC0FFFFFFFFFFFFFFFF0ABF0ABE0ABD0ABC0ABB0ABA0AB90AB8",
		x"0AD30AD20AD10AD00ACF0ACE0ACD0ACC0ACB0ACA0AC90AC80AC70AC60AC50AC4",
		x"0AE30AE20AE10AE00ADF0ADE0ADD0ADC0ADB0ADA0AD90AD80AD70AD60AD50AD4",
		x"0AF30AF20AF10AF00AEF0AEE0AED0AEC0AEB0AEA0AE90AE80AE70AE60AE50AE4",
		x"FFFFFFFFFFFFFFFF0AFF0AFE0AFD0AFC0AFB0AFA0AF90AF80AF70AF60AF50AF4",
		x"0B0F0B0E0B0D0B0C0B0B0B0A0B090B080B070B060B050B040B030B020B010B00",
		x"0B1F0B1E0B1D0B1C0B1B0B1A0B190B180B170B160B150B140B130B120B110B10",
		x"0B2F0B2E0B2D0B2C0B2B0B2A0B290B280B270B260B250B240B230B220B210B20",
		x"0B3F0B3E0B3D0B3C0B3B0B3A0B390B380B370B360B350B340B330B320B310B30",
		x"0B4B0B4A0B490B480B470B460B450B440B430B420B410B40FFFFFFFFFFFFFFFF",
		x"0B5B0B5A0B590B580B570B560B550B540B530B520B510B500B4F0B4E0B4D0B4C",
		x"0B6B0B6A0B690B680B670B660B650B640B630B620B610B600B5F0B5E0B5D0B5C",
		x"0B7B0B7A0B790B780B770B760B750B740B730B720B710B700B6F0B6E0B6D0B6C",
		x"0B870B860B850B840B830B820B810B80FFFFFFFFFFFFFFFF0B7F0B7E0B7D0B7C",
		x"0B970B960B950B940B930B920B910B900B8F0B8E0B8D0B8C0B8B0B8A0B890B88",
		x"0BA70BA60BA50BA40BA30BA20BA10BA00B9F0B9E0B9D0B9C0B9B0B9A0B990B98",
		x"0BB70BB60BB50BB40BB30BB20BB10BB00BAF0BAE0BAD0BAC0BAB0BAA0BA90BA8",
		x"0BC30BC20BC10BC0FFFFFFFFFFFFFFFF0BBF0BBE0BBD0BBC0BBB0BBA0BB90BB8",
		x"0BD30BD20BD10BD00BCF0BCE0BCD0BCC0BCB0BCA0BC90BC80BC70BC60BC50BC4",
		x"0BE30BE20BE10BE00BDF0BDE0BDD0BDC0BDB0BDA0BD90BD80BD70BD60BD50BD4",
		x"0BF30BF20BF10BF00BEF0BEE0BED0BEC0BEB0BEA0BE90BE80BE70BE60BE50BE4",
		x"FFFFFFFFFFFFFFFF0BFF0BFE0BFD0BFC0BFB0BFA0BF90BF80BF70BF60BF50BF4",
		x"0C0F0C0E0C0D0C0C0C0B0C0A0C090C080C070C060C050C040C030C020C010C00",
		x"0C1F0C1E0C1D0C1C0C1B0C1A0C190C180C170C160C150C140C130C120C110C10",
		x"0C2F0C2E0C2D0C2C0C2B0C2A0C290C280C270C260C250C240C230C220C210C20",
		x"0C3F0C3E0C3D0C3C0C3B0C3A0C390C380C370C360C350C340C330C320C310C30",
		x"0C4B0C4A0C490C480C470C460C450C440C430C420C410C40FFFFFFFFFFFFFFFF",
		x"0C5B0C5A0C590C580C570C560C550C540C530C520C510C500C4F0C4E0C4D0C4C",
		x"0C6B0C6A0C690C680C670C660C650C640C630C620C610C600C5F0C5E0C5D0C5C",
		x"0C7B0C7A0C790C780C770C760C750C740C730C720C710C700C6F0C6E0C6D0C6C",
		x"0C870C860C850C840C830C820C810C80FFFFFFFFFFFFFFFF0C7F0C7E0C7D0C7C",
		x"0C970C960C950C940C930C920C910C900C8F0C8E0C8D0C8C0C8B0C8A0C890C88",
		x"0CA70CA60CA50CA40CA30CA20CA10CA00C9F0C9E0C9D0C9C0C9B0C9A0C990C98",
		x"0CB70CB60CB50CB40CB30CB20CB10CB00CAF0CAE0CAD0CAC0CAB0CAA0CA90CA8",
		x"0CC30CC20CC10CC0FFFFFFFFFFFFFFFF0CBF0CBE0CBD0CBC0CBB0CBA0CB90CB8",
		x"0CD30CD20CD10CD00CCF0CCE0CCD0CCC0CCB0CCA0CC90CC80CC70CC60CC50CC4",
		x"0CE30CE20CE10CE00CDF0CDE0CDD0CDC0CDB0CDA0CD90CD80CD70CD60CD50CD4",
		x"0CF30CF20CF10CF00CEF0CEE0CED0CEC0CEB0CEA0CE90CE80CE70CE60CE50CE4",
		x"FFFFFFFFFFFFFFFF0CFF0CFE0CFD0CFC0CFB0CFA0CF90CF80CF70CF60CF50CF4",
		x"0D0F0D0E0D0D0D0C0D0B0D0A0D090D080D070D060D050D040D030D020D010D00",
		x"0D1F0D1E0D1D0D1C0D1B0D1A0D190D180D170D160D150D140D130D120D110D10",
		x"0D2F0D2E0D2D0D2C0D2B0D2A0D290D280D270D260D250D240D230D220D210D20",
		x"0D3F0D3E0D3D0D3C0D3B0D3A0D390D380D370D360D350D340D330D320D310D30",
		x"0D4B0D4A0D490D480D470D460D450D440D430D420D410D40FFFFFFFFFFFFFFFF",
		x"0D5B0D5A0D590D580D570D560D550D540D530D520D510D500D4F0D4E0D4D0D4C",
		x"0D6B0D6A0D690D680D670D660D650D640D630D620D610D600D5F0D5E0D5D0D5C",
		x"0D7B0D7A0D790D780D770D760D750D740D730D720D710D700D6F0D6E0D6D0D6C",
		x"0D870D860D850D840D830D820D810D80FFFFFFFFFFFFFFFF0D7F0D7E0D7D0D7C",
		x"0D970D960D950D940D930D920D910D900D8F0D8E0D8D0D8C0D8B0D8A0D890D88",
		x"0DA70DA60DA50DA40DA30DA20DA10DA00D9F0D9E0D9D0D9C0D9B0D9A0D990D98",
		x"0DB70DB60DB50DB40DB30DB20DB10DB00DAF0DAE0DAD0DAC0DAB0DAA0DA90DA8",
		x"0DC30DC20DC10DC0FFFFFFFFFFFFFFFF0DBF0DBE0DBD0DBC0DBB0DBA0DB90DB8",
		x"0DD30DD20DD10DD00DCF0DCE0DCD0DCC0DCB0DCA0DC90DC80DC70DC60DC50DC4",
		x"0DE30DE20DE10DE00DDF0DDE0DDD0DDC0DDB0DDA0DD90DD80DD70DD60DD50DD4",
		x"0DF30DF20DF10DF00DEF0DEE0DED0DEC0DEB0DEA0DE90DE80DE70DE60DE50DE4",
		x"FFFFFFFFFFFFFFFF0DFF0DFE0DFD0DFC0DFB0DFA0DF90DF80DF70DF60DF50DF4",
		x"0E0F0E0E0E0D0E0C0E0B0E0A0E090E080E070E060E050E040E030E020E010E00",
		x"0E1F0E1E0E1D0E1C0E1B0E1A0E190E180E170E160E150E140E130E120E110E10",
		x"0E2F0E2E0E2D0E2C0E2B0E2A0E290E280E270E260E250E240E230E220E210E20",
		x"0E3F0E3E0E3D0E3C0E3B0E3A0E390E380E370E360E350E340E330E320E310E30",
		x"0E4B0E4A0E490E480E470E460E450E440E430E420E410E40FFFFFFFFFFFFFFFF",
		x"0E5B0E5A0E590E580E570E560E550E540E530E520E510E500E4F0E4E0E4D0E4C",
		x"0E6B0E6A0E690E680E670E660E650E640E630E620E610E600E5F0E5E0E5D0E5C",
		x"0E7B0E7A0E790E780E770E760E750E740E730E720E710E700E6F0E6E0E6D0E6C",
		x"0E870E860E850E840E830E820E810E80FFFFFFFFFFFFFFFF0E7F0E7E0E7D0E7C",
		x"0E970E960E950E940E930E920E910E900E8F0E8E0E8D0E8C0E8B0E8A0E890E88",
		x"0EA70EA60EA50EA40EA30EA20EA10EA00E9F0E9E0E9D0E9C0E9B0E9A0E990E98",
		x"0EB70EB60EB50EB40EB30EB20EB10EB00EAF0EAE0EAD0EAC0EAB0EAA0EA90EA8",
		x"0EC30EC20EC10EC0FFFFFFFFFFFFFFFF0EBF0EBE0EBD0EBC0EBB0EBA0EB90EB8",
		x"0ED30ED20ED10ED00ECF0ECE0ECD0ECC0ECB0ECA0EC90EC80EC70EC60EC50EC4",
		x"0EE30EE20EE10EE00EDF0EDE0EDD0EDC0EDB0EDA0ED90ED80ED70ED60ED50ED4",
		x"0EF30EF20EF10EF00EEF0EEE0EED0EEC0EEB0EEA0EE90EE80EE70EE60EE50EE4",
		x"FFFFFFFFFFFFFFFF0EFF0EFE0EFD0EFC0EFB0EFA0EF90EF80EF70EF60EF50EF4",
		x"0F0F0F0E0F0D0F0C0F0B0F0A0F090F080F070F060F050F040F030F020F010F00",
		x"0F1F0F1E0F1D0F1C0F1B0F1A0F190F180F170F160F150F140F130F120F110F10",
		x"0F2F0F2E0F2D0F2C0F2B0F2A0F290F280F270F260F250F240F230F220F210F20",
		x"0F3F0F3E0F3D0F3C0F3B0F3A0F390F380F370F360F350F340F330F320F310F30",
		x"0F4B0F4A0F490F480F470F460F450F440F430F420F410F40FFFFFFFFFFFFFFFF",
		x"0F5B0F5A0F590F580F570F560F550F540F530F520F510F500F4F0F4E0F4D0F4C",
		x"0F6B0F6A0F690F680F670F660F650F640F630F620F610F600F5F0F5E0F5D0F5C",
		x"0F7B0F7A0F790F780F770F760F750F740F730F720F710F700F6F0F6E0F6D0F6C",
		x"0F870F860F850F840F830F820F810F80FFFFFFFFFFFFFFFF0F7F0F7E0F7D0F7C",
		x"0F970F960F950F940F930F920F910F900F8F0F8E0F8D0F8C0F8B0F8A0F890F88",
		x"0FA70FA60FA50FA40FA30FA20FA10FA00F9F0F9E0F9D0F9C0F9B0F9A0F990F98",
		x"0FB70FB60FB50FB40FB30FB20FB10FB00FAF0FAE0FAD0FAC0FAB0FAA0FA90FA8",
		x"0FC30FC20FC10FC0FFFFFFFFFFFFFFFF0FBF0FBE0FBD0FBC0FBB0FBA0FB90FB8",
		x"0FD30FD20FD10FD00FCF0FCE0FCD0FCC0FCB0FCA0FC90FC80FC70FC60FC50FC4",
		x"0FE30FE20FE10FE00FDF0FDE0FDD0FDC0FDB0FDA0FD90FD80FD70FD60FD50FD4",
		x"0FF30FF20FF10FF00FEF0FEE0FED0FEC0FEB0FEA0FE90FE80FE70FE60FE50FE4",
		x"FFFFFFFFFFFFFFFF0FFF0FFE0FFD0FFC0FFB0FFA0FF90FF80FF70FF60FF50FF4",
		x"100F100E100D100C100B100A1009100810071006100510041003100210011000",
		x"101F101E101D101C101B101A1019101810171016101510141013101210111010",
		x"102F102E102D102C102B102A1029102810271026102510241023102210211020",
		x"103F103E103D103C103B103A1039103810371036103510341033103210311030",
		x"104B104A1049104810471046104510441043104210411040FFFFFFFFFFFFFFFF",
		x"105B105A1059105810571056105510541053105210511050104F104E104D104C",
		x"106B106A1069106810671066106510641063106210611060105F105E105D105C",
		x"107B107A1079107810771076107510741073107210711070106F106E106D106C",
		x"10871086108510841083108210811080FFFFFFFFFFFFFFFF107F107E107D107C",
		x"10971096109510941093109210911090108F108E108D108C108B108A10891088",
		x"10A710A610A510A410A310A210A110A0109F109E109D109C109B109A10991098",
		x"10B710B610B510B410B310B210B110B010AF10AE10AD10AC10AB10AA10A910A8",
		x"10C310C210C110C0FFFFFFFFFFFFFFFF10BF10BE10BD10BC10BB10BA10B910B8",
		x"10D310D210D110D010CF10CE10CD10CC10CB10CA10C910C810C710C610C510C4",
		x"10E310E210E110E010DF10DE10DD10DC10DB10DA10D910D810D710D610D510D4",
		x"10F310F210F110F010EF10EE10ED10EC10EB10EA10E910E810E710E610E510E4",
		x"FFFFFFFFFFFFFFFF10FF10FE10FD10FC10FB10FA10F910F810F710F610F510F4",
		x"110F110E110D110C110B110A1109110811071106110511041103110211011100",
		x"111F111E111D111C111B111A1119111811171116111511141113111211111110",
		x"112F112E112D112C112B112A1129112811271126112511241123112211211120",
		x"113F113E113D113C113B113A1139113811371136113511341133113211311130",
		x"114B114A1149114811471146114511441143114211411140FFFFFFFFFFFFFFFF",
		x"115B115A1159115811571156115511541153115211511150114F114E114D114C",
		x"116B116A1169116811671166116511641163116211611160115F115E115D115C",
		x"117B117A1179117811771176117511741173117211711170116F116E116D116C",
		x"11871186118511841183118211811180FFFFFFFFFFFFFFFF117F117E117D117C",
		x"11971196119511941193119211911190118F118E118D118C118B118A11891188",
		x"11A711A611A511A411A311A211A111A0119F119E119D119C119B119A11991198",
		x"11B711B611B511B411B311B211B111B011AF11AE11AD11AC11AB11AA11A911A8",
		x"11C311C211C111C0FFFFFFFFFFFFFFFF11BF11BE11BD11BC11BB11BA11B911B8",
		x"11D311D211D111D011CF11CE11CD11CC11CB11CA11C911C811C711C611C511C4",
		x"11E311E211E111E011DF11DE11DD11DC11DB11DA11D911D811D711D611D511D4",
		x"11F311F211F111F011EF11EE11ED11EC11EB11EA11E911E811E711E611E511E4",
		x"FFFFFFFFFFFFFFFF11FF11FE11FD11FC11FB11FA11F911F811F711F611F511F4",
		x"120F120E120D120C120B120A1209120812071206120512041203120212011200",
		x"121F121E121D121C121B121A1219121812171216121512141213121212111210",
		x"122F122E122D122C122B122A1229122812271226122512241223122212211220",
		x"123F123E123D123C123B123A1239123812371236123512341233123212311230",
		x"124B124A1249124812471246124512441243124212411240FFFFFFFFFFFFFFFF",
		x"125B125A1259125812571256125512541253125212511250124F124E124D124C",
		x"126B126A1269126812671266126512641263126212611260125F125E125D125C",
		x"127B127A1279127812771276127512741273127212711270126F126E126D126C",
		x"12871286128512841283128212811280FFFFFFFFFFFFFFFF127F127E127D127C",
		x"12971296129512941293129212911290128F128E128D128C128B128A12891288",
		x"12A712A612A512A412A312A212A112A0129F129E129D129C129B129A12991298",
		x"12B712B612B512B412B312B212B112B012AF12AE12AD12AC12AB12AA12A912A8",
		x"12C312C212C112C0FFFFFFFFFFFFFFFF12BF12BE12BD12BC12BB12BA12B912B8",
		x"12D312D212D112D012CF12CE12CD12CC12CB12CA12C912C812C712C612C512C4",
		x"12E312E212E112E012DF12DE12DD12DC12DB12DA12D912D812D712D612D512D4",
		x"12F312F212F112F012EF12EE12ED12EC12EB12EA12E912E812E712E612E512E4",
		x"FFFFFFFFFFFFFFFF12FF12FE12FD12FC12FB12FA12F912F812F712F612F512F4",
		x"130F130E130D130C130B130A1309130813071306130513041303130213011300",
		x"131F131E131D131C131B131A1319131813171316131513141313131213111310",
		x"132F132E132D132C132B132A1329132813271326132513241323132213211320",
		x"133F133E133D133C133B133A1339133813371336133513341333133213311330",
		x"134B134A1349134813471346134513441343134213411340FFFFFFFFFFFFFFFF",
		x"135B135A1359135813571356135513541353135213511350134F134E134D134C",
		x"136B136A1369136813671366136513641363136213611360135F135E135D135C",
		x"137B137A1379137813771376137513741373137213711370136F136E136D136C",
		x"13871386138513841383138213811380FFFFFFFFFFFFFFFF137F137E137D137C",
		x"13971396139513941393139213911390138F138E138D138C138B138A13891388",
		x"13A713A613A513A413A313A213A113A0139F139E139D139C139B139A13991398",
		x"13B713B613B513B413B313B213B113B013AF13AE13AD13AC13AB13AA13A913A8",
		x"13C313C213C113C0FFFFFFFFFFFFFFFF13BF13BE13BD13BC13BB13BA13B913B8",
		x"13D313D213D113D013CF13CE13CD13CC13CB13CA13C913C813C713C613C513C4",
		x"13E313E213E113E013DF13DE13DD13DC13DB13DA13D913D813D713D613D513D4",
		x"13F313F213F113F013EF13EE13ED13EC13EB13EA13E913E813E713E613E513E4",
		x"FFFFFFFFFFFFFFFF13FF13FE13FD13FC13FB13FA13F913F813F713F613F513F4",
		x"140F140E140D140C140B140A1409140814071406140514041403140214011400",
		x"141F141E141D141C141B141A1419141814171416141514141413141214111410",
		x"142F142E142D142C142B142A1429142814271426142514241423142214211420",
		x"143F143E143D143C143B143A1439143814371436143514341433143214311430",
		x"144B144A1449144814471446144514441443144214411440FFFFFFFFFFFFFFFF",
		x"145B145A1459145814571456145514541453145214511450144F144E144D144C",
		x"146B146A1469146814671466146514641463146214611460145F145E145D145C",
		x"147B147A1479147814771476147514741473147214711470146F146E146D146C",
		x"14871486148514841483148214811480FFFFFFFFFFFFFFFF147F147E147D147C",
		x"14971496149514941493149214911490148F148E148D148C148B148A14891488",
		x"14A714A614A514A414A314A214A114A0149F149E149D149C149B149A14991498",
		x"14B714B614B514B414B314B214B114B014AF14AE14AD14AC14AB14AA14A914A8",
		x"14C314C214C114C0FFFFFFFFFFFFFFFF14BF14BE14BD14BC14BB14BA14B914B8",
		x"14D314D214D114D014CF14CE14CD14CC14CB14CA14C914C814C714C614C514C4",
		x"14E314E214E114E014DF14DE14DD14DC14DB14DA14D914D814D714D614D514D4",
		x"14F314F214F114F014EF14EE14ED14EC14EB14EA14E914E814E714E614E514E4",
		x"FFFFFFFFFFFFFFFF14FF14FE14FD14FC14FB14FA14F914F814F714F614F514F4",
		x"150F150E150D150C150B150A1509150815071506150515041503150215011500",
		x"151F151E151D151C151B151A1519151815171516151515141513151215111510",
		x"152F152E152D152C152B152A1529152815271526152515241523152215211520",
		x"153F153E153D153C153B153A1539153815371536153515341533153215311530",
		x"154B154A1549154815471546154515441543154215411540FFFFFFFFFFFFFFFF",
		x"155B155A1559155815571556155515541553155215511550154F154E154D154C",
		x"156B156A1569156815671566156515641563156215611560155F155E155D155C",
		x"157B157A1579157815771576157515741573157215711570156F156E156D156C",
		x"15871586158515841583158215811580FFFFFFFFFFFFFFFF157F157E157D157C",
		x"15971596159515941593159215911590158F158E158D158C158B158A15891588",
		x"15A715A615A515A415A315A215A115A0159F159E159D159C159B159A15991598",
		x"15B715B615B515B415B315B215B115B015AF15AE15AD15AC15AB15AA15A915A8",
		x"15C315C215C115C0FFFFFFFFFFFFFFFF15BF15BE15BD15BC15BB15BA15B915B8",
		x"15D315D215D115D015CF15CE15CD15CC15CB15CA15C915C815C715C615C515C4",
		x"15E315E215E115E015DF15DE15DD15DC15DB15DA15D915D815D715D615D515D4",
		x"15F315F215F115F015EF15EE15ED15EC15EB15EA15E915E815E715E615E515E4",
		x"FFFFFFFFFFFFFFFF15FF15FE15FD15FC15FB15FA15F915F815F715F615F515F4",
		x"160F160E160D160C160B160A1609160816071606160516041603160216011600",
		x"161F161E161D161C161B161A1619161816171616161516141613161216111610",
		x"162F162E162D162C162B162A1629162816271626162516241623162216211620",
		x"163F163E163D163C163B163A1639163816371636163516341633163216311630",
		x"164B164A1649164816471646164516441643164216411640FFFFFFFFFFFFFFFF",
		x"165B165A1659165816571656165516541653165216511650164F164E164D164C",
		x"166B166A1669166816671666166516641663166216611660165F165E165D165C",
		x"167B167A1679167816771676167516741673167216711670166F166E166D166C",
		x"16871686168516841683168216811680FFFFFFFFFFFFFFFF167F167E167D167C",
		x"16971696169516941693169216911690168F168E168D168C168B168A16891688",
		x"16A716A616A516A416A316A216A116A0169F169E169D169C169B169A16991698",
		x"16B716B616B516B416B316B216B116B016AF16AE16AD16AC16AB16AA16A916A8",
		x"16C316C216C116C0FFFFFFFFFFFFFFFF16BF16BE16BD16BC16BB16BA16B916B8",
		x"16D316D216D116D016CF16CE16CD16CC16CB16CA16C916C816C716C616C516C4",
		x"16E316E216E116E016DF16DE16DD16DC16DB16DA16D916D816D716D616D516D4",
		x"16F316F216F116F016EF16EE16ED16EC16EB16EA16E916E816E716E616E516E4",
		x"FFFFFFFFFFFFFFFF16FF16FE16FD16FC16FB16FA16F916F816F716F616F516F4",
		x"170F170E170D170C170B170A1709170817071706170517041703170217011700",
		x"171F171E171D171C171B171A1719171817171716171517141713171217111710",
		x"172F172E172D172C172B172A1729172817271726172517241723172217211720",
		x"173F173E173D173C173B173A1739173817371736173517341733173217311730",
		x"174B174A1749174817471746174517441743174217411740FFFFFFFFFFFFFFFF",
		x"175B175A1759175817571756175517541753175217511750174F174E174D174C",
		x"176B176A1769176817671766176517641763176217611760175F175E175D175C",
		x"177B177A1779177817771776177517741773177217711770176F176E176D176C",
		x"17871786178517841783178217811780FFFFFFFFFFFFFFFF177F177E177D177C",
		x"17971796179517941793179217911790178F178E178D178C178B178A17891788",
		x"17A717A617A517A417A317A217A117A0179F179E179D179C179B179A17991798",
		x"17B717B617B517B417B317B217B117B017AF17AE17AD17AC17AB17AA17A917A8",
		x"17C317C217C117C0FFFFFFFFFFFFFFFF17BF17BE17BD17BC17BB17BA17B917B8",
		x"17D317D217D117D017CF17CE17CD17CC17CB17CA17C917C817C717C617C517C4",
		x"17E317E217E117E017DF17DE17DD17DC17DB17DA17D917D817D717D617D517D4",
		x"17F317F217F117F017EF17EE17ED17EC17EB17EA17E917E817E717E617E517E4",
		x"FFFFFFFFFFFFFFFF17FF17FE17FD17FC17FB17FA17F917F817F717F617F517F4",
		x"180F180E180D180C180B180A1809180818071806180518041803180218011800",
		x"181F181E181D181C181B181A1819181818171816181518141813181218111810",
		x"182F182E182D182C182B182A1829182818271826182518241823182218211820",
		x"183F183E183D183C183B183A1839183818371836183518341833183218311830",
		x"184B184A1849184818471846184518441843184218411840FFFFFFFFFFFFFFFF",
		x"185B185A1859185818571856185518541853185218511850184F184E184D184C",
		x"186B186A1869186818671866186518641863186218611860185F185E185D185C",
		x"187B187A1879187818771876187518741873187218711870186F186E186D186C",
		x"18871886188518841883188218811880FFFFFFFFFFFFFFFF187F187E187D187C",
		x"18971896189518941893189218911890188F188E188D188C188B188A18891888",
		x"18A718A618A518A418A318A218A118A0189F189E189D189C189B189A18991898",
		x"18B718B618B518B418B318B218B118B018AF18AE18AD18AC18AB18AA18A918A8",
		x"18C318C218C118C0FFFFFFFFFFFFFFFF18BF18BE18BD18BC18BB18BA18B918B8",
		x"18D318D218D118D018CF18CE18CD18CC18CB18CA18C918C818C718C618C518C4",
		x"18E318E218E118E018DF18DE18DD18DC18DB18DA18D918D818D718D618D518D4",
		x"18F318F218F118F018EF18EE18ED18EC18EB18EA18E918E818E718E618E518E4",
		x"FFFFFFFFFFFFFFFF18FF18FE18FD18FC18FB18FA18F918F818F718F618F518F4",
		x"190F190E190D190C190B190A1909190819071906190519041903190219011900",
		x"191F191E191D191C191B191A1919191819171916191519141913191219111910",
		x"192F192E192D192C192B192A1929192819271926192519241923192219211920",
		x"193F193E193D193C193B193A1939193819371936193519341933193219311930",
		x"194B194A1949194819471946194519441943194219411940FFFFFFFFFFFFFFFF",
		x"195B195A1959195819571956195519541953195219511950194F194E194D194C",
		x"196B196A1969196819671966196519641963196219611960195F195E195D195C",
		x"197B197A1979197819771976197519741973197219711970196F196E196D196C",
		x"19871986198519841983198219811980FFFFFFFFFFFFFFFF197F197E197D197C",
		x"19971996199519941993199219911990198F198E198D198C198B198A19891988",
		x"19A719A619A519A419A319A219A119A0199F199E199D199C199B199A19991998",
		x"19B719B619B519B419B319B219B119B019AF19AE19AD19AC19AB19AA19A919A8",
		x"19C319C219C119C0FFFFFFFFFFFFFFFF19BF19BE19BD19BC19BB19BA19B919B8",
		x"19D319D219D119D019CF19CE19CD19CC19CB19CA19C919C819C719C619C519C4",
		x"19E319E219E119E019DF19DE19DD19DC19DB19DA19D919D819D719D619D519D4",
		x"19F319F219F119F019EF19EE19ED19EC19EB19EA19E919E819E719E619E519E4",
		x"FFFFFFFFFFFFFFFF19FF19FE19FD19FC19FB19FA19F919F819F719F619F519F4",
		x"1A0F1A0E1A0D1A0C1A0B1A0A1A091A081A071A061A051A041A031A021A011A00",
		x"1A1F1A1E1A1D1A1C1A1B1A1A1A191A181A171A161A151A141A131A121A111A10",
		x"1A2F1A2E1A2D1A2C1A2B1A2A1A291A281A271A261A251A241A231A221A211A20",
		x"1A3F1A3E1A3D1A3C1A3B1A3A1A391A381A371A361A351A341A331A321A311A30",
		x"1A4B1A4A1A491A481A471A461A451A441A431A421A411A40FFFFFFFFFFFFFFFF",
		x"1A5B1A5A1A591A581A571A561A551A541A531A521A511A501A4F1A4E1A4D1A4C",
		x"1A6B1A6A1A691A681A671A661A651A641A631A621A611A601A5F1A5E1A5D1A5C",
		x"1A7B1A7A1A791A781A771A761A751A741A731A721A711A701A6F1A6E1A6D1A6C",
		x"1A871A861A851A841A831A821A811A80FFFFFFFFFFFFFFFF1A7F1A7E1A7D1A7C",
		x"1A971A961A951A941A931A921A911A901A8F1A8E1A8D1A8C1A8B1A8A1A891A88",
		x"1AA71AA61AA51AA41AA31AA21AA11AA01A9F1A9E1A9D1A9C1A9B1A9A1A991A98",
		x"1AB71AB61AB51AB41AB31AB21AB11AB01AAF1AAE1AAD1AAC1AAB1AAA1AA91AA8",
		x"1AC31AC21AC11AC0FFFFFFFFFFFFFFFF1ABF1ABE1ABD1ABC1ABB1ABA1AB91AB8",
		x"1AD31AD21AD11AD01ACF1ACE1ACD1ACC1ACB1ACA1AC91AC81AC71AC61AC51AC4",
		x"1AE31AE21AE11AE01ADF1ADE1ADD1ADC1ADB1ADA1AD91AD81AD71AD61AD51AD4",
		x"1AF31AF21AF11AF01AEF1AEE1AED1AEC1AEB1AEA1AE91AE81AE71AE61AE51AE4",
		x"FFFFFFFFFFFFFFFF1AFF1AFE1AFD1AFC1AFB1AFA1AF91AF81AF71AF61AF51AF4",
		x"1B0F1B0E1B0D1B0C1B0B1B0A1B091B081B071B061B051B041B031B021B011B00",
		x"1B1F1B1E1B1D1B1C1B1B1B1A1B191B181B171B161B151B141B131B121B111B10",
		x"1B2F1B2E1B2D1B2C1B2B1B2A1B291B281B271B261B251B241B231B221B211B20",
		x"1B3F1B3E1B3D1B3C1B3B1B3A1B391B381B371B361B351B341B331B321B311B30",
		x"1B4B1B4A1B491B481B471B461B451B441B431B421B411B40FFFFFFFFFFFFFFFF",
		x"1B5B1B5A1B591B581B571B561B551B541B531B521B511B501B4F1B4E1B4D1B4C",
		x"1B6B1B6A1B691B681B671B661B651B641B631B621B611B601B5F1B5E1B5D1B5C",
		x"1B7B1B7A1B791B781B771B761B751B741B731B721B711B701B6F1B6E1B6D1B6C",
		x"1B871B861B851B841B831B821B811B80FFFFFFFFFFFFFFFF1B7F1B7E1B7D1B7C",
		x"1B971B961B951B941B931B921B911B901B8F1B8E1B8D1B8C1B8B1B8A1B891B88",
		x"1BA71BA61BA51BA41BA31BA21BA11BA01B9F1B9E1B9D1B9C1B9B1B9A1B991B98",
		x"1BB71BB61BB51BB41BB31BB21BB11BB01BAF1BAE1BAD1BAC1BAB1BAA1BA91BA8",
		x"1BC31BC21BC11BC0FFFFFFFFFFFFFFFF1BBF1BBE1BBD1BBC1BBB1BBA1BB91BB8",
		x"1BD31BD21BD11BD01BCF1BCE1BCD1BCC1BCB1BCA1BC91BC81BC71BC61BC51BC4",
		x"1BE31BE21BE11BE01BDF1BDE1BDD1BDC1BDB1BDA1BD91BD81BD71BD61BD51BD4",
		x"1BF31BF21BF11BF01BEF1BEE1BED1BEC1BEB1BEA1BE91BE81BE71BE61BE51BE4",
		x"FFFFFFFFFFFFFFFF1BFF1BFE1BFD1BFC1BFB1BFA1BF91BF81BF71BF61BF51BF4",
		x"1C0F1C0E1C0D1C0C1C0B1C0A1C091C081C071C061C051C041C031C021C011C00",
		x"1C1F1C1E1C1D1C1C1C1B1C1A1C191C181C171C161C151C141C131C121C111C10",
		x"1C2F1C2E1C2D1C2C1C2B1C2A1C291C281C271C261C251C241C231C221C211C20",
		x"1C3F1C3E1C3D1C3C1C3B1C3A1C391C381C371C361C351C341C331C321C311C30",
		x"1C4B1C4A1C491C481C471C461C451C441C431C421C411C40FFFFFFFFFFFFFFFF",
		x"1C5B1C5A1C591C581C571C561C551C541C531C521C511C501C4F1C4E1C4D1C4C",
		x"1C6B1C6A1C691C681C671C661C651C641C631C621C611C601C5F1C5E1C5D1C5C",
		x"1C7B1C7A1C791C781C771C761C751C741C731C721C711C701C6F1C6E1C6D1C6C",
		x"1C871C861C851C841C831C821C811C80FFFFFFFFFFFFFFFF1C7F1C7E1C7D1C7C",
		x"1C971C961C951C941C931C921C911C901C8F1C8E1C8D1C8C1C8B1C8A1C891C88",
		x"1CA71CA61CA51CA41CA31CA21CA11CA01C9F1C9E1C9D1C9C1C9B1C9A1C991C98",
		x"1CB71CB61CB51CB41CB31CB21CB11CB01CAF1CAE1CAD1CAC1CAB1CAA1CA91CA8",
		x"1CC31CC21CC11CC0FFFFFFFFFFFFFFFF1CBF1CBE1CBD1CBC1CBB1CBA1CB91CB8",
		x"1CD31CD21CD11CD01CCF1CCE1CCD1CCC1CCB1CCA1CC91CC81CC71CC61CC51CC4",
		x"1CE31CE21CE11CE01CDF1CDE1CDD1CDC1CDB1CDA1CD91CD81CD71CD61CD51CD4",
		x"1CF31CF21CF11CF01CEF1CEE1CED1CEC1CEB1CEA1CE91CE81CE71CE61CE51CE4",
		x"FFFFFFFFFFFFFFFF1CFF1CFE1CFD1CFC1CFB1CFA1CF91CF81CF71CF61CF51CF4",
		x"1D0F1D0E1D0D1D0C1D0B1D0A1D091D081D071D061D051D041D031D021D011D00",
		x"1D1F1D1E1D1D1D1C1D1B1D1A1D191D181D171D161D151D141D131D121D111D10",
		x"1D2F1D2E1D2D1D2C1D2B1D2A1D291D281D271D261D251D241D231D221D211D20",
		x"1D3F1D3E1D3D1D3C1D3B1D3A1D391D381D371D361D351D341D331D321D311D30",
		x"1D4B1D4A1D491D481D471D461D451D441D431D421D411D40FFFFFFFFFFFFFFFF",
		x"1D5B1D5A1D591D581D571D561D551D541D531D521D511D501D4F1D4E1D4D1D4C",
		x"1D6B1D6A1D691D681D671D661D651D641D631D621D611D601D5F1D5E1D5D1D5C",
		x"1D7B1D7A1D791D781D771D761D751D741D731D721D711D701D6F1D6E1D6D1D6C",
		x"1D871D861D851D841D831D821D811D80FFFFFFFFFFFFFFFF1D7F1D7E1D7D1D7C",
		x"1D971D961D951D941D931D921D911D901D8F1D8E1D8D1D8C1D8B1D8A1D891D88",
		x"1DA71DA61DA51DA41DA31DA21DA11DA01D9F1D9E1D9D1D9C1D9B1D9A1D991D98",
		x"1DB71DB61DB51DB41DB31DB21DB11DB01DAF1DAE1DAD1DAC1DAB1DAA1DA91DA8",
		x"1DC31DC21DC11DC0FFFFFFFFFFFFFFFF1DBF1DBE1DBD1DBC1DBB1DBA1DB91DB8",
		x"1DD31DD21DD11DD01DCF1DCE1DCD1DCC1DCB1DCA1DC91DC81DC71DC61DC51DC4",
		x"1DE31DE21DE11DE01DDF1DDE1DDD1DDC1DDB1DDA1DD91DD81DD71DD61DD51DD4",
		x"1DF31DF21DF11DF01DEF1DEE1DED1DEC1DEB1DEA1DE91DE81DE71DE61DE51DE4",
		x"FFFFFFFFFFFFFFFF1DFF1DFE1DFD1DFC1DFB1DFA1DF91DF81DF71DF61DF51DF4",
		x"1E0F1E0E1E0D1E0C1E0B1E0A1E091E081E071E061E051E041E031E021E011E00",
		x"1E1F1E1E1E1D1E1C1E1B1E1A1E191E181E171E161E151E141E131E121E111E10",
		x"1E2F1E2E1E2D1E2C1E2B1E2A1E291E281E271E261E251E241E231E221E211E20",
		x"1E3F1E3E1E3D1E3C1E3B1E3A1E391E381E371E361E351E341E331E321E311E30",
		x"1E4B1E4A1E491E481E471E461E451E441E431E421E411E40FFFFFFFFFFFFFFFF",
		x"1E5B1E5A1E591E581E571E561E551E541E531E521E511E501E4F1E4E1E4D1E4C",
		x"1E6B1E6A1E691E681E671E661E651E641E631E621E611E601E5F1E5E1E5D1E5C",
		x"1E7B1E7A1E791E781E771E761E751E741E731E721E711E701E6F1E6E1E6D1E6C",
		x"1E871E861E851E841E831E821E811E80FFFFFFFFFFFFFFFF1E7F1E7E1E7D1E7C",
		x"1E971E961E951E941E931E921E911E901E8F1E8E1E8D1E8C1E8B1E8A1E891E88",
		x"1EA71EA61EA51EA41EA31EA21EA11EA01E9F1E9E1E9D1E9C1E9B1E9A1E991E98",
		x"1EB71EB61EB51EB41EB31EB21EB11EB01EAF1EAE1EAD1EAC1EAB1EAA1EA91EA8",
		x"1EC31EC21EC11EC0FFFFFFFFFFFFFFFF1EBF1EBE1EBD1EBC1EBB1EBA1EB91EB8",
		x"1ED31ED21ED11ED01ECF1ECE1ECD1ECC1ECB1ECA1EC91EC81EC71EC61EC51EC4",
		x"1EE31EE21EE11EE01EDF1EDE1EDD1EDC1EDB1EDA1ED91ED81ED71ED61ED51ED4",
		x"1EF31EF21EF11EF01EEF1EEE1EED1EEC1EEB1EEA1EE91EE81EE71EE61EE51EE4",
		x"FFFFFFFFFFFFFFFF1EFF1EFE1EFD1EFC1EFB1EFA1EF91EF81EF71EF61EF51EF4",
		x"1F0F1F0E1F0D1F0C1F0B1F0A1F091F081F071F061F051F041F031F021F011F00",
		x"1F1F1F1E1F1D1F1C1F1B1F1A1F191F181F171F161F151F141F131F121F111F10",
		x"1F2F1F2E1F2D1F2C1F2B1F2A1F291F281F271F261F251F241F231F221F211F20",
		x"1F3F1F3E1F3D1F3C1F3B1F3A1F391F381F371F361F351F341F331F321F311F30",
		x"1F4B1F4A1F491F481F471F461F451F441F431F421F411F40FFFFFFFFFFFFFFFF",
		x"1F5B1F5A1F591F581F571F561F551F541F531F521F511F501F4F1F4E1F4D1F4C",
		x"1F6B1F6A1F691F681F671F661F651F641F631F621F611F601F5F1F5E1F5D1F5C",
		x"1F7B1F7A1F791F781F771F761F751F741F731F721F711F701F6F1F6E1F6D1F6C",
		x"1F871F861F851F841F831F821F811F80FFFFFFFFFFFFFFFF1F7F1F7E1F7D1F7C",
		x"1F971F961F951F941F931F921F911F901F8F1F8E1F8D1F8C1F8B1F8A1F891F88",
		x"1FA71FA61FA51FA41FA31FA21FA11FA01F9F1F9E1F9D1F9C1F9B1F9A1F991F98",
		x"1FB71FB61FB51FB41FB31FB21FB11FB01FAF1FAE1FAD1FAC1FAB1FAA1FA91FA8",
		x"1FC31FC21FC11FC0FFFFFFFFFFFFFFFF1FBF1FBE1FBD1FBC1FBB1FBA1FB91FB8",
		x"1FD31FD21FD11FD01FCF1FCE1FCD1FCC1FCB1FCA1FC91FC81FC71FC61FC51FC4",
		x"1FE31FE21FE11FE01FDF1FDE1FDD1FDC1FDB1FDA1FD91FD81FD71FD61FD51FD4",
		x"1FF31FF21FF11FF01FEF1FEE1FED1FEC1FEB1FEA1FE91FE81FE71FE61FE51FE4",
		x"FFFFFFFFFFFFFFFF1FFF1FFE1FFD1FFC1FFB1FFA1FF91FF81FF71FF61FF51FF4",
		x"200F200E200D200C200B200A2009200820072006200520042003200220012000",
		x"201F201E201D201C201B201A2019201820172016201520142013201220112010",
		x"202F202E202D202C202B202A2029202820272026202520242023202220212020",
		x"203F203E203D203C203B203A2039203820372036203520342033203220312030",
		x"204B204A2049204820472046204520442043204220412040FFFFFFFFFFFFFFFF",
		x"205B205A2059205820572056205520542053205220512050204F204E204D204C",
		x"206B206A2069206820672066206520642063206220612060205F205E205D205C",
		x"207B207A2079207820772076207520742073207220712070206F206E206D206C",
		x"20872086208520842083208220812080FFFFFFFFFFFFFFFF207F207E207D207C",
		x"20972096209520942093209220912090208F208E208D208C208B208A20892088",
		x"20A720A620A520A420A320A220A120A0209F209E209D209C209B209A20992098",
		x"20B720B620B520B420B320B220B120B020AF20AE20AD20AC20AB20AA20A920A8",
		x"20C320C220C120C0FFFFFFFFFFFFFFFF20BF20BE20BD20BC20BB20BA20B920B8",
		x"20D320D220D120D020CF20CE20CD20CC20CB20CA20C920C820C720C620C520C4",
		x"20E320E220E120E020DF20DE20DD20DC20DB20DA20D920D820D720D620D520D4",
		x"20F320F220F120F020EF20EE20ED20EC20EB20EA20E920E820E720E620E520E4",
		x"FFFFFFFFFFFFFFFF20FF20FE20FD20FC20FB20FA20F920F820F720F620F520F4",
		x"210F210E210D210C210B210A2109210821072106210521042103210221012100",
		x"211F211E211D211C211B211A2119211821172116211521142113211221112110",
		x"212F212E212D212C212B212A2129212821272126212521242123212221212120",
		x"213F213E213D213C213B213A2139213821372136213521342133213221312130",
		x"214B214A2149214821472146214521442143214221412140FFFFFFFFFFFFFFFF",
		x"215B215A2159215821572156215521542153215221512150214F214E214D214C",
		x"216B216A2169216821672166216521642163216221612160215F215E215D215C",
		x"217B217A2179217821772176217521742173217221712170216F216E216D216C",
		x"21872186218521842183218221812180FFFFFFFFFFFFFFFF217F217E217D217C",
		x"21972196219521942193219221912190218F218E218D218C218B218A21892188",
		x"21A721A621A521A421A321A221A121A0219F219E219D219C219B219A21992198",
		x"21B721B621B521B421B321B221B121B021AF21AE21AD21AC21AB21AA21A921A8",
		x"21C321C221C121C0FFFFFFFFFFFFFFFF21BF21BE21BD21BC21BB21BA21B921B8",
		x"21D321D221D121D021CF21CE21CD21CC21CB21CA21C921C821C721C621C521C4",
		x"21E321E221E121E021DF21DE21DD21DC21DB21DA21D921D821D721D621D521D4",
		x"21F321F221F121F021EF21EE21ED21EC21EB21EA21E921E821E721E621E521E4",
		x"FFFFFFFFFFFFFFFF21FF21FE21FD21FC21FB21FA21F921F821F721F621F521F4",
		x"220F220E220D220C220B220A2209220822072206220522042203220222012200",
		x"221F221E221D221C221B221A2219221822172216221522142213221222112210",
		x"222F222E222D222C222B222A2229222822272226222522242223222222212220",
		x"223F223E223D223C223B223A2239223822372236223522342233223222312230",
		x"224B224A2249224822472246224522442243224222412240FFFFFFFFFFFFFFFF",
		x"225B225A2259225822572256225522542253225222512250224F224E224D224C",
		x"226B226A2269226822672266226522642263226222612260225F225E225D225C",
		x"227B227A2279227822772276227522742273227222712270226F226E226D226C",
		x"22872286228522842283228222812280FFFFFFFFFFFFFFFF227F227E227D227C",
		x"22972296229522942293229222912290228F228E228D228C228B228A22892288",
		x"22A722A622A522A422A322A222A122A0229F229E229D229C229B229A22992298",
		x"22B722B622B522B422B322B222B122B022AF22AE22AD22AC22AB22AA22A922A8",
		x"22C322C222C122C0FFFFFFFFFFFFFFFF22BF22BE22BD22BC22BB22BA22B922B8",
		x"22D322D222D122D022CF22CE22CD22CC22CB22CA22C922C822C722C622C522C4",
		x"22E322E222E122E022DF22DE22DD22DC22DB22DA22D922D822D722D622D522D4",
		x"22F322F222F122F022EF22EE22ED22EC22EB22EA22E922E822E722E622E522E4",
		x"FFFFFFFFFFFFFFFF22FF22FE22FD22FC22FB22FA22F922F822F722F622F522F4",
		x"230F230E230D230C230B230A2309230823072306230523042303230223012300",
		x"231F231E231D231C231B231A2319231823172316231523142313231223112310",
		x"232F232E232D232C232B232A2329232823272326232523242323232223212320",
		x"233F233E233D233C233B233A2339233823372336233523342333233223312330",
		x"234B234A2349234823472346234523442343234223412340FFFFFFFFFFFFFFFF",
		x"235B235A2359235823572356235523542353235223512350234F234E234D234C",
		x"236B236A2369236823672366236523642363236223612360235F235E235D235C",
		x"237B237A2379237823772376237523742373237223712370236F236E236D236C",
		x"23872386238523842383238223812380FFFFFFFFFFFFFFFF237F237E237D237C",
		x"23972396239523942393239223912390238F238E238D238C238B238A23892388",
		x"23A723A623A523A423A323A223A123A0239F239E239D239C239B239A23992398",
		x"23B723B623B523B423B323B223B123B023AF23AE23AD23AC23AB23AA23A923A8",
		x"23C323C223C123C0FFFFFFFFFFFFFFFF23BF23BE23BD23BC23BB23BA23B923B8",
		x"23D323D223D123D023CF23CE23CD23CC23CB23CA23C923C823C723C623C523C4",
		x"23E323E223E123E023DF23DE23DD23DC23DB23DA23D923D823D723D623D523D4",
		x"23F323F223F123F023EF23EE23ED23EC23EB23EA23E923E823E723E623E523E4",
		x"FFFFFFFFFFFFFFFF23FF23FE23FD23FC23FB23FA23F923F823F723F623F523F4",
		x"240F240E240D240C240B240A2409240824072406240524042403240224012400",
		x"241F241E241D241C241B241A2419241824172416241524142413241224112410",
		x"242F242E242D242C242B242A2429242824272426242524242423242224212420",
		x"243F243E243D243C243B243A2439243824372436243524342433243224312430",
		x"244B244A2449244824472446244524442443244224412440FFFFFFFFFFFFFFFF",
		x"245B245A2459245824572456245524542453245224512450244F244E244D244C",
		x"246B246A2469246824672466246524642463246224612460245F245E245D245C",
		x"247B247A2479247824772476247524742473247224712470246F246E246D246C",
		x"24872486248524842483248224812480FFFFFFFFFFFFFFFF247F247E247D247C",
		x"24972496249524942493249224912490248F248E248D248C248B248A24892488",
		x"24A724A624A524A424A324A224A124A0249F249E249D249C249B249A24992498",
		x"24B724B624B524B424B324B224B124B024AF24AE24AD24AC24AB24AA24A924A8",
		x"24C324C224C124C0FFFFFFFFFFFFFFFF24BF24BE24BD24BC24BB24BA24B924B8",
		x"24D324D224D124D024CF24CE24CD24CC24CB24CA24C924C824C724C624C524C4",
		x"24E324E224E124E024DF24DE24DD24DC24DB24DA24D924D824D724D624D524D4",
		x"24F324F224F124F024EF24EE24ED24EC24EB24EA24E924E824E724E624E524E4",
		x"FFFFFFFFFFFFFFFF24FF24FE24FD24FC24FB24FA24F924F824F724F624F524F4",
		x"250F250E250D250C250B250A2509250825072506250525042503250225012500",
		x"251F251E251D251C251B251A2519251825172516251525142513251225112510",
		x"252F252E252D252C252B252A2529252825272526252525242523252225212520",
		x"253F253E253D253C253B253A2539253825372536253525342533253225312530",
		x"254B254A2549254825472546254525442543254225412540FFFFFFFFFFFFFFFF",
		x"255B255A2559255825572556255525542553255225512550254F254E254D254C",
		x"256B256A2569256825672566256525642563256225612560255F255E255D255C",
		x"257B257A2579257825772576257525742573257225712570256F256E256D256C",
		x"25872586258525842583258225812580FFFFFFFFFFFFFFFF257F257E257D257C",
		x"25972596259525942593259225912590258F258E258D258C258B258A25892588",
		x"25A725A625A525A425A325A225A125A0259F259E259D259C259B259A25992598",
		x"25B725B625B525B425B325B225B125B025AF25AE25AD25AC25AB25AA25A925A8",
		x"25C325C225C125C0FFFFFFFFFFFFFFFF25BF25BE25BD25BC25BB25BA25B925B8",
		x"25D325D225D125D025CF25CE25CD25CC25CB25CA25C925C825C725C625C525C4",
		x"25E325E225E125E025DF25DE25DD25DC25DB25DA25D925D825D725D625D525D4",
		x"25F325F225F125F025EF25EE25ED25EC25EB25EA25E925E825E725E625E525E4",
		x"FFFFFFFFFFFFFFFF25FF25FE25FD25FC25FB25FA25F925F825F725F625F525F4",
		x"260F260E260D260C260B260A2609260826072606260526042603260226012600",
		x"261F261E261D261C261B261A2619261826172616261526142613261226112610",
		x"262F262E262D262C262B262A2629262826272626262526242623262226212620",
		x"263F263E263D263C263B263A2639263826372636263526342633263226312630",
		x"264B264A2649264826472646264526442643264226412640FFFFFFFFFFFFFFFF",
		x"265B265A2659265826572656265526542653265226512650264F264E264D264C",
		x"266B266A2669266826672666266526642663266226612660265F265E265D265C",
		x"267B267A2679267826772676267526742673267226712670266F266E266D266C",
		x"26872686268526842683268226812680FFFFFFFFFFFFFFFF267F267E267D267C",
		x"26972696269526942693269226912690268F268E268D268C268B268A26892688",
		x"26A726A626A526A426A326A226A126A0269F269E269D269C269B269A26992698",
		x"26B726B626B526B426B326B226B126B026AF26AE26AD26AC26AB26AA26A926A8",
		x"26C326C226C126C0FFFFFFFFFFFFFFFF26BF26BE26BD26BC26BB26BA26B926B8",
		x"26D326D226D126D026CF26CE26CD26CC26CB26CA26C926C826C726C626C526C4",
		x"26E326E226E126E026DF26DE26DD26DC26DB26DA26D926D826D726D626D526D4",
		x"26F326F226F126F026EF26EE26ED26EC26EB26EA26E926E826E726E626E526E4",
		x"FFFFFFFFFFFFFFFF26FF26FE26FD26FC26FB26FA26F926F826F726F626F526F4",
		x"270F270E270D270C270B270A2709270827072706270527042703270227012700",
		x"271F271E271D271C271B271A2719271827172716271527142713271227112710",
		x"272F272E272D272C272B272A2729272827272726272527242723272227212720",
		x"273F273E273D273C273B273A2739273827372736273527342733273227312730",
		x"274B274A2749274827472746274527442743274227412740FFFFFFFFFFFFFFFF",
		x"275B275A2759275827572756275527542753275227512750274F274E274D274C",
		x"276B276A2769276827672766276527642763276227612760275F275E275D275C",
		x"277B277A2779277827772776277527742773277227712770276F276E276D276C",
		x"27872786278527842783278227812780FFFFFFFFFFFFFFFF277F277E277D277C",
		x"27972796279527942793279227912790278F278E278D278C278B278A27892788",
		x"27A727A627A527A427A327A227A127A0279F279E279D279C279B279A27992798",
		x"27B727B627B527B427B327B227B127B027AF27AE27AD27AC27AB27AA27A927A8",
		x"27C327C227C127C0FFFFFFFFFFFFFFFF27BF27BE27BD27BC27BB27BA27B927B8",
		x"27D327D227D127D027CF27CE27CD27CC27CB27CA27C927C827C727C627C527C4",
		x"27E327E227E127E027DF27DE27DD27DC27DB27DA27D927D827D727D627D527D4",
		x"27F327F227F127F027EF27EE27ED27EC27EB27EA27E927E827E727E627E527E4",
		x"FFFFFFFFFFFFFFFF27FF27FE27FD27FC27FB27FA27F927F827F727F627F527F4",
		x"280F280E280D280C280B280A2809280828072806280528042803280228012800",
		x"281F281E281D281C281B281A2819281828172816281528142813281228112810",
		x"282F282E282D282C282B282A2829282828272826282528242823282228212820",
		x"283F283E283D283C283B283A2839283828372836283528342833283228312830",
		x"284B284A2849284828472846284528442843284228412840FFFFFFFFFFFFFFFF",
		x"285B285A2859285828572856285528542853285228512850284F284E284D284C",
		x"286B286A2869286828672866286528642863286228612860285F285E285D285C",
		x"287B287A2879287828772876287528742873287228712870286F286E286D286C",
		x"28872886288528842883288228812880FFFFFFFFFFFFFFFF287F287E287D287C",
		x"28972896289528942893289228912890288F288E288D288C288B288A28892888",
		x"28A728A628A528A428A328A228A128A0289F289E289D289C289B289A28992898",
		x"28B728B628B528B428B328B228B128B028AF28AE28AD28AC28AB28AA28A928A8",
		x"28C328C228C128C0FFFFFFFFFFFFFFFF28BF28BE28BD28BC28BB28BA28B928B8",
		x"28D328D228D128D028CF28CE28CD28CC28CB28CA28C928C828C728C628C528C4",
		x"28E328E228E128E028DF28DE28DD28DC28DB28DA28D928D828D728D628D528D4",
		x"28F328F228F128F028EF28EE28ED28EC28EB28EA28E928E828E728E628E528E4",
		x"FFFFFFFFFFFFFFFF28FF28FE28FD28FC28FB28FA28F928F828F728F628F528F4",
		x"290F290E290D290C290B290A2909290829072906290529042903290229012900",
		x"291F291E291D291C291B291A2919291829172916291529142913291229112910",
		x"292F292E292D292C292B292A2929292829272926292529242923292229212920",
		x"293F293E293D293C293B293A2939293829372936293529342933293229312930",
		x"294B294A2949294829472946294529442943294229412940FFFFFFFFFFFFFFFF",
		x"295B295A2959295829572956295529542953295229512950294F294E294D294C",
		x"296B296A2969296829672966296529642963296229612960295F295E295D295C",
		x"297B297A2979297829772976297529742973297229712970296F296E296D296C",
		x"29872986298529842983298229812980FFFFFFFFFFFFFFFF297F297E297D297C",
		x"29972996299529942993299229912990298F298E298D298C298B298A29892988",
		x"29A729A629A529A429A329A229A129A0299F299E299D299C299B299A29992998",
		x"29B729B629B529B429B329B229B129B029AF29AE29AD29AC29AB29AA29A929A8",
		x"29C329C229C129C0FFFFFFFFFFFFFFFF29BF29BE29BD29BC29BB29BA29B929B8",
		x"29D329D229D129D029CF29CE29CD29CC29CB29CA29C929C829C729C629C529C4",
		x"29E329E229E129E029DF29DE29DD29DC29DB29DA29D929D829D729D629D529D4",
		x"29F329F229F129F029EF29EE29ED29EC29EB29EA29E929E829E729E629E529E4",
		x"FFFFFFFFFFFFFFFF29FF29FE29FD29FC29FB29FA29F929F829F729F629F529F4",
		x"2A0F2A0E2A0D2A0C2A0B2A0A2A092A082A072A062A052A042A032A022A012A00",
		x"2A1F2A1E2A1D2A1C2A1B2A1A2A192A182A172A162A152A142A132A122A112A10",
		x"2A2F2A2E2A2D2A2C2A2B2A2A2A292A282A272A262A252A242A232A222A212A20",
		x"2A3F2A3E2A3D2A3C2A3B2A3A2A392A382A372A362A352A342A332A322A312A30",
		x"2A4B2A4A2A492A482A472A462A452A442A432A422A412A40FFFFFFFFFFFFFFFF",
		x"2A5B2A5A2A592A582A572A562A552A542A532A522A512A502A4F2A4E2A4D2A4C",
		x"2A6B2A6A2A692A682A672A662A652A642A632A622A612A602A5F2A5E2A5D2A5C",
		x"2A7B2A7A2A792A782A772A762A752A742A732A722A712A702A6F2A6E2A6D2A6C",
		x"2A872A862A852A842A832A822A812A80FFFFFFFFFFFFFFFF2A7F2A7E2A7D2A7C",
		x"2A972A962A952A942A932A922A912A902A8F2A8E2A8D2A8C2A8B2A8A2A892A88",
		x"2AA72AA62AA52AA42AA32AA22AA12AA02A9F2A9E2A9D2A9C2A9B2A9A2A992A98",
		x"2AB72AB62AB52AB42AB32AB22AB12AB02AAF2AAE2AAD2AAC2AAB2AAA2AA92AA8",
		x"2AC32AC22AC12AC0FFFFFFFFFFFFFFFF2ABF2ABE2ABD2ABC2ABB2ABA2AB92AB8",
		x"2AD32AD22AD12AD02ACF2ACE2ACD2ACC2ACB2ACA2AC92AC82AC72AC62AC52AC4",
		x"2AE32AE22AE12AE02ADF2ADE2ADD2ADC2ADB2ADA2AD92AD82AD72AD62AD52AD4",
		x"2AF32AF22AF12AF02AEF2AEE2AED2AEC2AEB2AEA2AE92AE82AE72AE62AE52AE4",
		x"FFFFFFFFFFFFFFFF2AFF2AFE2AFD2AFC2AFB2AFA2AF92AF82AF72AF62AF52AF4",
		x"2B0F2B0E2B0D2B0C2B0B2B0A2B092B082B072B062B052B042B032B022B012B00",
		x"2B1F2B1E2B1D2B1C2B1B2B1A2B192B182B172B162B152B142B132B122B112B10",
		x"2B2F2B2E2B2D2B2C2B2B2B2A2B292B282B272B262B252B242B232B222B212B20",
		x"2B3F2B3E2B3D2B3C2B3B2B3A2B392B382B372B362B352B342B332B322B312B30",
		x"2B4B2B4A2B492B482B472B462B452B442B432B422B412B40FFFFFFFFFFFFFFFF",
		x"2B5B2B5A2B592B582B572B562B552B542B532B522B512B502B4F2B4E2B4D2B4C",
		x"2B6B2B6A2B692B682B672B662B652B642B632B622B612B602B5F2B5E2B5D2B5C",
		x"2B7B2B7A2B792B782B772B762B752B742B732B722B712B702B6F2B6E2B6D2B6C",
		x"2B872B862B852B842B832B822B812B80FFFFFFFFFFFFFFFF2B7F2B7E2B7D2B7C",
		x"2B972B962B952B942B932B922B912B902B8F2B8E2B8D2B8C2B8B2B8A2B892B88",
		x"2BA72BA62BA52BA42BA32BA22BA12BA02B9F2B9E2B9D2B9C2B9B2B9A2B992B98",
		x"2BB72BB62BB52BB42BB32BB22BB12BB02BAF2BAE2BAD2BAC2BAB2BAA2BA92BA8",
		x"2BC32BC22BC12BC0FFFFFFFFFFFFFFFF2BBF2BBE2BBD2BBC2BBB2BBA2BB92BB8",
		x"2BD32BD22BD12BD02BCF2BCE2BCD2BCC2BCB2BCA2BC92BC82BC72BC62BC52BC4",
		x"2BE32BE22BE12BE02BDF2BDE2BDD2BDC2BDB2BDA2BD92BD82BD72BD62BD52BD4",
		x"2BF32BF22BF12BF02BEF2BEE2BED2BEC2BEB2BEA2BE92BE82BE72BE62BE52BE4",
		x"FFFFFFFFFFFFFFFF2BFF2BFE2BFD2BFC2BFB2BFA2BF92BF82BF72BF62BF52BF4",
		x"2C0F2C0E2C0D2C0C2C0B2C0A2C092C082C072C062C052C042C032C022C012C00",
		x"2C1F2C1E2C1D2C1C2C1B2C1A2C192C182C172C162C152C142C132C122C112C10",
		x"2C2F2C2E2C2D2C2C2C2B2C2A2C292C282C272C262C252C242C232C222C212C20",
		x"2C3F2C3E2C3D2C3C2C3B2C3A2C392C382C372C362C352C342C332C322C312C30",
		x"2C4B2C4A2C492C482C472C462C452C442C432C422C412C40FFFFFFFFFFFFFFFF",
		x"2C5B2C5A2C592C582C572C562C552C542C532C522C512C502C4F2C4E2C4D2C4C",
		x"2C6B2C6A2C692C682C672C662C652C642C632C622C612C602C5F2C5E2C5D2C5C",
		x"2C7B2C7A2C792C782C772C762C752C742C732C722C712C702C6F2C6E2C6D2C6C",
		x"2C872C862C852C842C832C822C812C80FFFFFFFFFFFFFFFF2C7F2C7E2C7D2C7C",
		x"2C972C962C952C942C932C922C912C902C8F2C8E2C8D2C8C2C8B2C8A2C892C88",
		x"2CA72CA62CA52CA42CA32CA22CA12CA02C9F2C9E2C9D2C9C2C9B2C9A2C992C98",
		x"2CB72CB62CB52CB42CB32CB22CB12CB02CAF2CAE2CAD2CAC2CAB2CAA2CA92CA8",
		x"2CC32CC22CC12CC0FFFFFFFFFFFFFFFF2CBF2CBE2CBD2CBC2CBB2CBA2CB92CB8",
		x"2CD32CD22CD12CD02CCF2CCE2CCD2CCC2CCB2CCA2CC92CC82CC72CC62CC52CC4",
		x"2CE32CE22CE12CE02CDF2CDE2CDD2CDC2CDB2CDA2CD92CD82CD72CD62CD52CD4",
		x"2CF32CF22CF12CF02CEF2CEE2CED2CEC2CEB2CEA2CE92CE82CE72CE62CE52CE4",
		x"FFFFFFFFFFFFFFFF2CFF2CFE2CFD2CFC2CFB2CFA2CF92CF82CF72CF62CF52CF4",
		x"2D0F2D0E2D0D2D0C2D0B2D0A2D092D082D072D062D052D042D032D022D012D00",
		x"2D1F2D1E2D1D2D1C2D1B2D1A2D192D182D172D162D152D142D132D122D112D10",
		x"2D2F2D2E2D2D2D2C2D2B2D2A2D292D282D272D262D252D242D232D222D212D20",
		x"2D3F2D3E2D3D2D3C2D3B2D3A2D392D382D372D362D352D342D332D322D312D30",
		x"2D4B2D4A2D492D482D472D462D452D442D432D422D412D40FFFFFFFFFFFFFFFF",
		x"2D5B2D5A2D592D582D572D562D552D542D532D522D512D502D4F2D4E2D4D2D4C",
		x"2D6B2D6A2D692D682D672D662D652D642D632D622D612D602D5F2D5E2D5D2D5C",
		x"2D7B2D7A2D792D782D772D762D752D742D732D722D712D702D6F2D6E2D6D2D6C",
		x"2D872D862D852D842D832D822D812D80FFFFFFFFFFFFFFFF2D7F2D7E2D7D2D7C",
		x"2D972D962D952D942D932D922D912D902D8F2D8E2D8D2D8C2D8B2D8A2D892D88",
		x"2DA72DA62DA52DA42DA32DA22DA12DA02D9F2D9E2D9D2D9C2D9B2D9A2D992D98",
		x"2DB72DB62DB52DB42DB32DB22DB12DB02DAF2DAE2DAD2DAC2DAB2DAA2DA92DA8",
		x"2DC32DC22DC12DC0FFFFFFFFFFFFFFFF2DBF2DBE2DBD2DBC2DBB2DBA2DB92DB8",
		x"2DD32DD22DD12DD02DCF2DCE2DCD2DCC2DCB2DCA2DC92DC82DC72DC62DC52DC4",
		x"2DE32DE22DE12DE02DDF2DDE2DDD2DDC2DDB2DDA2DD92DD82DD72DD62DD52DD4",
		x"2DF32DF22DF12DF02DEF2DEE2DED2DEC2DEB2DEA2DE92DE82DE72DE62DE52DE4",
		x"FFFFFFFFFFFFFFFF2DFF2DFE2DFD2DFC2DFB2DFA2DF92DF82DF72DF62DF52DF4",
		x"2E0F2E0E2E0D2E0C2E0B2E0A2E092E082E072E062E052E042E032E022E012E00",
		x"2E1F2E1E2E1D2E1C2E1B2E1A2E192E182E172E162E152E142E132E122E112E10",
		x"2E2F2E2E2E2D2E2C2E2B2E2A2E292E282E272E262E252E242E232E222E212E20",
		x"2E3F2E3E2E3D2E3C2E3B2E3A2E392E382E372E362E352E342E332E322E312E30",
		x"2E4B2E4A2E492E482E472E462E452E442E432E422E412E40FFFFFFFFFFFFFFFF",
		x"2E5B2E5A2E592E582E572E562E552E542E532E522E512E502E4F2E4E2E4D2E4C",
		x"2E6B2E6A2E692E682E672E662E652E642E632E622E612E602E5F2E5E2E5D2E5C",
		x"2E7B2E7A2E792E782E772E762E752E742E732E722E712E702E6F2E6E2E6D2E6C",
		x"2E872E862E852E842E832E822E812E80FFFFFFFFFFFFFFFF2E7F2E7E2E7D2E7C",
		x"2E972E962E952E942E932E922E912E902E8F2E8E2E8D2E8C2E8B2E8A2E892E88",
		x"2EA72EA62EA52EA42EA32EA22EA12EA02E9F2E9E2E9D2E9C2E9B2E9A2E992E98",
		x"2EB72EB62EB52EB42EB32EB22EB12EB02EAF2EAE2EAD2EAC2EAB2EAA2EA92EA8",
		x"2EC32EC22EC12EC0FFFFFFFFFFFFFFFF2EBF2EBE2EBD2EBC2EBB2EBA2EB92EB8",
		x"2ED32ED22ED12ED02ECF2ECE2ECD2ECC2ECB2ECA2EC92EC82EC72EC62EC52EC4",
		x"2EE32EE22EE12EE02EDF2EDE2EDD2EDC2EDB2EDA2ED92ED82ED72ED62ED52ED4",
		x"2EF32EF22EF12EF02EEF2EEE2EED2EEC2EEB2EEA2EE92EE82EE72EE62EE52EE4",
		x"FFFFFFFFFFFFFFFF2EFF2EFE2EFD2EFC2EFB2EFA2EF92EF82EF72EF62EF52EF4",
		x"2F0F2F0E2F0D2F0C2F0B2F0A2F092F082F072F062F052F042F032F022F012F00",
		x"2F1F2F1E2F1D2F1C2F1B2F1A2F192F182F172F162F152F142F132F122F112F10",
		x"2F2F2F2E2F2D2F2C2F2B2F2A2F292F282F272F262F252F242F232F222F212F20",
		x"2F3F2F3E2F3D2F3C2F3B2F3A2F392F382F372F362F352F342F332F322F312F30",
		x"2F4B2F4A2F492F482F472F462F452F442F432F422F412F40FFFFFFFFFFFFFFFF",
		x"2F5B2F5A2F592F582F572F562F552F542F532F522F512F502F4F2F4E2F4D2F4C",
		x"2F6B2F6A2F692F682F672F662F652F642F632F622F612F602F5F2F5E2F5D2F5C",
		x"2F7B2F7A2F792F782F772F762F752F742F732F722F712F702F6F2F6E2F6D2F6C",
		x"2F872F862F852F842F832F822F812F80FFFFFFFFFFFFFFFF2F7F2F7E2F7D2F7C",
		x"2F972F962F952F942F932F922F912F902F8F2F8E2F8D2F8C2F8B2F8A2F892F88",
		x"2FA72FA62FA52FA42FA32FA22FA12FA02F9F2F9E2F9D2F9C2F9B2F9A2F992F98",
		x"2FB72FB62FB52FB42FB32FB22FB12FB02FAF2FAE2FAD2FAC2FAB2FAA2FA92FA8",
		x"2FC32FC22FC12FC0FFFFFFFFFFFFFFFF2FBF2FBE2FBD2FBC2FBB2FBA2FB92FB8",
		x"2FD32FD22FD12FD02FCF2FCE2FCD2FCC2FCB2FCA2FC92FC82FC72FC62FC52FC4",
		x"2FE32FE22FE12FE02FDF2FDE2FDD2FDC2FDB2FDA2FD92FD82FD72FD62FD52FD4",
		x"2FF32FF22FF12FF02FEF2FEE2FED2FEC2FEB2FEA2FE92FE82FE72FE62FE52FE4",
		x"FFFFFFFFFFFFFFFF2FFF2FFE2FFD2FFC2FFB2FFA2FF92FF82FF72FF62FF52FF4",
		x"300F300E300D300C300B300A3009300830073006300530043003300230013000",
		x"301F301E301D301C301B301A3019301830173016301530143013301230113010",
		x"302F302E302D302C302B302A3029302830273026302530243023302230213020",
		x"303F303E303D303C303B303A3039303830373036303530343033303230313030",
		x"304B304A3049304830473046304530443043304230413040FFFFFFFFFFFFFFFF",
		x"305B305A3059305830573056305530543053305230513050304F304E304D304C",
		x"306B306A3069306830673066306530643063306230613060305F305E305D305C",
		x"307B307A3079307830773076307530743073307230713070306F306E306D306C",
		x"30873086308530843083308230813080FFFFFFFFFFFFFFFF307F307E307D307C",
		x"30973096309530943093309230913090308F308E308D308C308B308A30893088",
		x"30A730A630A530A430A330A230A130A0309F309E309D309C309B309A30993098",
		x"30B730B630B530B430B330B230B130B030AF30AE30AD30AC30AB30AA30A930A8",
		x"30C330C230C130C0FFFFFFFFFFFFFFFF30BF30BE30BD30BC30BB30BA30B930B8",
		x"30D330D230D130D030CF30CE30CD30CC30CB30CA30C930C830C730C630C530C4",
		x"30E330E230E130E030DF30DE30DD30DC30DB30DA30D930D830D730D630D530D4",
		x"30F330F230F130F030EF30EE30ED30EC30EB30EA30E930E830E730E630E530E4",
		x"FFFFFFFFFFFFFFFF30FF30FE30FD30FC30FB30FA30F930F830F730F630F530F4",
		x"310F310E310D310C310B310A3109310831073106310531043103310231013100",
		x"311F311E311D311C311B311A3119311831173116311531143113311231113110",
		x"312F312E312D312C312B312A3129312831273126312531243123312231213120",
		x"313F313E313D313C313B313A3139313831373136313531343133313231313130",
		x"314B314A3149314831473146314531443143314231413140FFFFFFFFFFFFFFFF",
		x"315B315A3159315831573156315531543153315231513150314F314E314D314C",
		x"316B316A3169316831673166316531643163316231613160315F315E315D315C",
		x"317B317A3179317831773176317531743173317231713170316F316E316D316C",
		x"31873186318531843183318231813180FFFFFFFFFFFFFFFF317F317E317D317C",
		x"31973196319531943193319231913190318F318E318D318C318B318A31893188",
		x"31A731A631A531A431A331A231A131A0319F319E319D319C319B319A31993198",
		x"31B731B631B531B431B331B231B131B031AF31AE31AD31AC31AB31AA31A931A8",
		x"31C331C231C131C0FFFFFFFFFFFFFFFF31BF31BE31BD31BC31BB31BA31B931B8",
		x"31D331D231D131D031CF31CE31CD31CC31CB31CA31C931C831C731C631C531C4",
		x"31E331E231E131E031DF31DE31DD31DC31DB31DA31D931D831D731D631D531D4",
		x"31F331F231F131F031EF31EE31ED31EC31EB31EA31E931E831E731E631E531E4",
		x"FFFFFFFFFFFFFFFF31FF31FE31FD31FC31FB31FA31F931F831F731F631F531F4",
		x"320F320E320D320C320B320A3209320832073206320532043203320232013200",
		x"321F321E321D321C321B321A3219321832173216321532143213321232113210",
		x"322F322E322D322C322B322A3229322832273226322532243223322232213220",
		x"323F323E323D323C323B323A3239323832373236323532343233323232313230",
		x"324B324A3249324832473246324532443243324232413240FFFFFFFFFFFFFFFF",
		x"325B325A3259325832573256325532543253325232513250324F324E324D324C",
		x"326B326A3269326832673266326532643263326232613260325F325E325D325C",
		x"327B327A3279327832773276327532743273327232713270326F326E326D326C",
		x"32873286328532843283328232813280FFFFFFFFFFFFFFFF327F327E327D327C",
		x"32973296329532943293329232913290328F328E328D328C328B328A32893288",
		x"32A732A632A532A432A332A232A132A0329F329E329D329C329B329A32993298",
		x"32B732B632B532B432B332B232B132B032AF32AE32AD32AC32AB32AA32A932A8",
		x"32C332C232C132C0FFFFFFFFFFFFFFFF32BF32BE32BD32BC32BB32BA32B932B8",
		x"32D332D232D132D032CF32CE32CD32CC32CB32CA32C932C832C732C632C532C4",
		x"32E332E232E132E032DF32DE32DD32DC32DB32DA32D932D832D732D632D532D4",
		x"32F332F232F132F032EF32EE32ED32EC32EB32EA32E932E832E732E632E532E4",
		x"FFFFFFFFFFFFFFFF32FF32FE32FD32FC32FB32FA32F932F832F732F632F532F4",
		x"330F330E330D330C330B330A3309330833073306330533043303330233013300",
		x"331F331E331D331C331B331A3319331833173316331533143313331233113310",
		x"332F332E332D332C332B332A3329332833273326332533243323332233213320",
		x"333F333E333D333C333B333A3339333833373336333533343333333233313330",
		x"334B334A3349334833473346334533443343334233413340FFFFFFFFFFFFFFFF",
		x"335B335A3359335833573356335533543353335233513350334F334E334D334C",
		x"336B336A3369336833673366336533643363336233613360335F335E335D335C",
		x"337B337A3379337833773376337533743373337233713370336F336E336D336C",
		x"33873386338533843383338233813380FFFFFFFFFFFFFFFF337F337E337D337C",
		x"33973396339533943393339233913390338F338E338D338C338B338A33893388",
		x"33A733A633A533A433A333A233A133A0339F339E339D339C339B339A33993398",
		x"33B733B633B533B433B333B233B133B033AF33AE33AD33AC33AB33AA33A933A8",
		x"33C333C233C133C0FFFFFFFFFFFFFFFF33BF33BE33BD33BC33BB33BA33B933B8",
		x"33D333D233D133D033CF33CE33CD33CC33CB33CA33C933C833C733C633C533C4",
		x"33E333E233E133E033DF33DE33DD33DC33DB33DA33D933D833D733D633D533D4",
		x"33F333F233F133F033EF33EE33ED33EC33EB33EA33E933E833E733E633E533E4",
		x"FFFFFFFFFFFFFFFF33FF33FE33FD33FC33FB33FA33F933F833F733F633F533F4",
		x"340F340E340D340C340B340A3409340834073406340534043403340234013400",
		x"341F341E341D341C341B341A3419341834173416341534143413341234113410",
		x"342F342E342D342C342B342A3429342834273426342534243423342234213420",
		x"343F343E343D343C343B343A3439343834373436343534343433343234313430",
		x"344B344A3449344834473446344534443443344234413440FFFFFFFFFFFFFFFF",
		x"345B345A3459345834573456345534543453345234513450344F344E344D344C",
		x"346B346A3469346834673466346534643463346234613460345F345E345D345C",
		x"347B347A3479347834773476347534743473347234713470346F346E346D346C",
		x"34873486348534843483348234813480FFFFFFFFFFFFFFFF347F347E347D347C",
		x"34973496349534943493349234913490348F348E348D348C348B348A34893488",
		x"34A734A634A534A434A334A234A134A0349F349E349D349C349B349A34993498",
		x"34B734B634B534B434B334B234B134B034AF34AE34AD34AC34AB34AA34A934A8",
		x"34C334C234C134C0FFFFFFFFFFFFFFFF34BF34BE34BD34BC34BB34BA34B934B8",
		x"34D334D234D134D034CF34CE34CD34CC34CB34CA34C934C834C734C634C534C4",
		x"34E334E234E134E034DF34DE34DD34DC34DB34DA34D934D834D734D634D534D4",
		x"34F334F234F134F034EF34EE34ED34EC34EB34EA34E934E834E734E634E534E4",
		x"FFFFFFFFFFFFFFFF34FF34FE34FD34FC34FB34FA34F934F834F734F634F534F4",
		x"350F350E350D350C350B350A3509350835073506350535043503350235013500",
		x"351F351E351D351C351B351A3519351835173516351535143513351235113510",
		x"352F352E352D352C352B352A3529352835273526352535243523352235213520",
		x"353F353E353D353C353B353A3539353835373536353535343533353235313530",
		x"354B354A3549354835473546354535443543354235413540FFFFFFFFFFFFFFFF",
		x"355B355A3559355835573556355535543553355235513550354F354E354D354C",
		x"356B356A3569356835673566356535643563356235613560355F355E355D355C",
		x"357B357A3579357835773576357535743573357235713570356F356E356D356C",
		x"35873586358535843583358235813580FFFFFFFFFFFFFFFF357F357E357D357C",
		x"35973596359535943593359235913590358F358E358D358C358B358A35893588",
		x"35A735A635A535A435A335A235A135A0359F359E359D359C359B359A35993598",
		x"35B735B635B535B435B335B235B135B035AF35AE35AD35AC35AB35AA35A935A8",
		x"35C335C235C135C0FFFFFFFFFFFFFFFF35BF35BE35BD35BC35BB35BA35B935B8",
		x"35D335D235D135D035CF35CE35CD35CC35CB35CA35C935C835C735C635C535C4",
		x"35E335E235E135E035DF35DE35DD35DC35DB35DA35D935D835D735D635D535D4",
		x"35F335F235F135F035EF35EE35ED35EC35EB35EA35E935E835E735E635E535E4",
		x"FFFFFFFFFFFFFFFF35FF35FE35FD35FC35FB35FA35F935F835F735F635F535F4",
		x"360F360E360D360C360B360A3609360836073606360536043603360236013600",
		x"361F361E361D361C361B361A3619361836173616361536143613361236113610",
		x"362F362E362D362C362B362A3629362836273626362536243623362236213620",
		x"363F363E363D363C363B363A3639363836373636363536343633363236313630",
		x"364B364A3649364836473646364536443643364236413640FFFFFFFFFFFFFFFF",
		x"365B365A3659365836573656365536543653365236513650364F364E364D364C",
		x"366B366A3669366836673666366536643663366236613660365F365E365D365C",
		x"367B367A3679367836773676367536743673367236713670366F366E366D366C",
		x"36873686368536843683368236813680FFFFFFFFFFFFFFFF367F367E367D367C",
		x"36973696369536943693369236913690368F368E368D368C368B368A36893688",
		x"36A736A636A536A436A336A236A136A0369F369E369D369C369B369A36993698",
		x"36B736B636B536B436B336B236B136B036AF36AE36AD36AC36AB36AA36A936A8",
		x"36C336C236C136C0FFFFFFFFFFFFFFFF36BF36BE36BD36BC36BB36BA36B936B8",
		x"36D336D236D136D036CF36CE36CD36CC36CB36CA36C936C836C736C636C536C4",
		x"36E336E236E136E036DF36DE36DD36DC36DB36DA36D936D836D736D636D536D4",
		x"36F336F236F136F036EF36EE36ED36EC36EB36EA36E936E836E736E636E536E4",
		x"FFFFFFFFFFFFFFFF36FF36FE36FD36FC36FB36FA36F936F836F736F636F536F4",
		x"370F370E370D370C370B370A3709370837073706370537043703370237013700",
		x"371F371E371D371C371B371A3719371837173716371537143713371237113710",
		x"372F372E372D372C372B372A3729372837273726372537243723372237213720",
		x"373F373E373D373C373B373A3739373837373736373537343733373237313730",
		x"374B374A3749374837473746374537443743374237413740FFFFFFFFFFFFFFFF",
		x"375B375A3759375837573756375537543753375237513750374F374E374D374C",
		x"376B376A3769376837673766376537643763376237613760375F375E375D375C",
		x"377B377A3779377837773776377537743773377237713770376F376E376D376C",
		x"37873786378537843783378237813780FFFFFFFFFFFFFFFF377F377E377D377C",
		x"37973796379537943793379237913790378F378E378D378C378B378A37893788",
		x"37A737A637A537A437A337A237A137A0379F379E379D379C379B379A37993798",
		x"37B737B637B537B437B337B237B137B037AF37AE37AD37AC37AB37AA37A937A8",
		x"37C337C237C137C0FFFFFFFFFFFFFFFF37BF37BE37BD37BC37BB37BA37B937B8",
		x"37D337D237D137D037CF37CE37CD37CC37CB37CA37C937C837C737C637C537C4",
		x"37E337E237E137E037DF37DE37DD37DC37DB37DA37D937D837D737D637D537D4",
		x"37F337F237F137F037EF37EE37ED37EC37EB37EA37E937E837E737E637E537E4",
		x"FFFFFFFFFFFFFFFF37FF37FE37FD37FC37FB37FA37F937F837F737F637F537F4",
		x"380F380E380D380C380B380A3809380838073806380538043803380238013800",
		x"381F381E381D381C381B381A3819381838173816381538143813381238113810",
		x"382F382E382D382C382B382A3829382838273826382538243823382238213820",
		x"383F383E383D383C383B383A3839383838373836383538343833383238313830",
		x"384B384A3849384838473846384538443843384238413840FFFFFFFFFFFFFFFF",
		x"385B385A3859385838573856385538543853385238513850384F384E384D384C",
		x"386B386A3869386838673866386538643863386238613860385F385E385D385C",
		x"387B387A3879387838773876387538743873387238713870386F386E386D386C",
		x"38873886388538843883388238813880FFFFFFFFFFFFFFFF387F387E387D387C",
		x"38973896389538943893389238913890388F388E388D388C388B388A38893888",
		x"38A738A638A538A438A338A238A138A0389F389E389D389C389B389A38993898",
		x"38B738B638B538B438B338B238B138B038AF38AE38AD38AC38AB38AA38A938A8",
		x"38C338C238C138C0FFFFFFFFFFFFFFFF38BF38BE38BD38BC38BB38BA38B938B8",
		x"38D338D238D138D038CF38CE38CD38CC38CB38CA38C938C838C738C638C538C4",
		x"38E338E238E138E038DF38DE38DD38DC38DB38DA38D938D838D738D638D538D4",
		x"38F338F238F138F038EF38EE38ED38EC38EB38EA38E938E838E738E638E538E4",
		x"FFFFFFFFFFFFFFFF38FF38FE38FD38FC38FB38FA38F938F838F738F638F538F4",
		x"390F390E390D390C390B390A3909390839073906390539043903390239013900",
		x"391F391E391D391C391B391A3919391839173916391539143913391239113910",
		x"392F392E392D392C392B392A3929392839273926392539243923392239213920",
		x"393F393E393D393C393B393A3939393839373936393539343933393239313930",
		x"394B394A3949394839473946394539443943394239413940FFFFFFFFFFFFFFFF",
		x"395B395A3959395839573956395539543953395239513950394F394E394D394C",
		x"396B396A3969396839673966396539643963396239613960395F395E395D395C",
		x"397B397A3979397839773976397539743973397239713970396F396E396D396C",
		x"39873986398539843983398239813980FFFFFFFFFFFFFFFF397F397E397D397C",
		x"39973996399539943993399239913990398F398E398D398C398B398A39893988",
		x"39A739A639A539A439A339A239A139A0399F399E399D399C399B399A39993998",
		x"39B739B639B539B439B339B239B139B039AF39AE39AD39AC39AB39AA39A939A8",
		x"39C339C239C139C0FFFFFFFFFFFFFFFF39BF39BE39BD39BC39BB39BA39B939B8",
		x"39D339D239D139D039CF39CE39CD39CC39CB39CA39C939C839C739C639C539C4",
		x"39E339E239E139E039DF39DE39DD39DC39DB39DA39D939D839D739D639D539D4",
		x"39F339F239F139F039EF39EE39ED39EC39EB39EA39E939E839E739E639E539E4",
		x"FFFFFFFFFFFFFFFF39FF39FE39FD39FC39FB39FA39F939F839F739F639F539F4",
		x"3A0F3A0E3A0D3A0C3A0B3A0A3A093A083A073A063A053A043A033A023A013A00",
		x"3A1F3A1E3A1D3A1C3A1B3A1A3A193A183A173A163A153A143A133A123A113A10",
		x"3A2F3A2E3A2D3A2C3A2B3A2A3A293A283A273A263A253A243A233A223A213A20",
		x"3A3F3A3E3A3D3A3C3A3B3A3A3A393A383A373A363A353A343A333A323A313A30",
		x"3A4B3A4A3A493A483A473A463A453A443A433A423A413A40FFFFFFFFFFFFFFFF",
		x"3A5B3A5A3A593A583A573A563A553A543A533A523A513A503A4F3A4E3A4D3A4C",
		x"3A6B3A6A3A693A683A673A663A653A643A633A623A613A603A5F3A5E3A5D3A5C",
		x"3A7B3A7A3A793A783A773A763A753A743A733A723A713A703A6F3A6E3A6D3A6C",
		x"3A873A863A853A843A833A823A813A80FFFFFFFFFFFFFFFF3A7F3A7E3A7D3A7C",
		x"3A973A963A953A943A933A923A913A903A8F3A8E3A8D3A8C3A8B3A8A3A893A88",
		x"3AA73AA63AA53AA43AA33AA23AA13AA03A9F3A9E3A9D3A9C3A9B3A9A3A993A98",
		x"3AB73AB63AB53AB43AB33AB23AB13AB03AAF3AAE3AAD3AAC3AAB3AAA3AA93AA8",
		x"3AC33AC23AC13AC0FFFFFFFFFFFFFFFF3ABF3ABE3ABD3ABC3ABB3ABA3AB93AB8",
		x"3AD33AD23AD13AD03ACF3ACE3ACD3ACC3ACB3ACA3AC93AC83AC73AC63AC53AC4",
		x"3AE33AE23AE13AE03ADF3ADE3ADD3ADC3ADB3ADA3AD93AD83AD73AD63AD53AD4",
		x"3AF33AF23AF13AF03AEF3AEE3AED3AEC3AEB3AEA3AE93AE83AE73AE63AE53AE4",
		x"FFFFFFFFFFFFFFFF3AFF3AFE3AFD3AFC3AFB3AFA3AF93AF83AF73AF63AF53AF4",
		x"3B0F3B0E3B0D3B0C3B0B3B0A3B093B083B073B063B053B043B033B023B013B00",
		x"3B1F3B1E3B1D3B1C3B1B3B1A3B193B183B173B163B153B143B133B123B113B10",
		x"3B2F3B2E3B2D3B2C3B2B3B2A3B293B283B273B263B253B243B233B223B213B20",
		x"3B3F3B3E3B3D3B3C3B3B3B3A3B393B383B373B363B353B343B333B323B313B30",
		x"3B4B3B4A3B493B483B473B463B453B443B433B423B413B40FFFFFFFFFFFFFFFF",
		x"3B5B3B5A3B593B583B573B563B553B543B533B523B513B503B4F3B4E3B4D3B4C",
		x"3B6B3B6A3B693B683B673B663B653B643B633B623B613B603B5F3B5E3B5D3B5C",
		x"3B7B3B7A3B793B783B773B763B753B743B733B723B713B703B6F3B6E3B6D3B6C",
		x"3B873B863B853B843B833B823B813B80FFFFFFFFFFFFFFFF3B7F3B7E3B7D3B7C",
		x"3B973B963B953B943B933B923B913B903B8F3B8E3B8D3B8C3B8B3B8A3B893B88",
		x"3BA73BA63BA53BA43BA33BA23BA13BA03B9F3B9E3B9D3B9C3B9B3B9A3B993B98",
		x"3BB73BB63BB53BB43BB33BB23BB13BB03BAF3BAE3BAD3BAC3BAB3BAA3BA93BA8",
		x"3BC33BC23BC13BC0FFFFFFFFFFFFFFFF3BBF3BBE3BBD3BBC3BBB3BBA3BB93BB8",
		x"3BD33BD23BD13BD03BCF3BCE3BCD3BCC3BCB3BCA3BC93BC83BC73BC63BC53BC4",
		x"3BE33BE23BE13BE03BDF3BDE3BDD3BDC3BDB3BDA3BD93BD83BD73BD63BD53BD4",
		x"3BF33BF23BF13BF03BEF3BEE3BED3BEC3BEB3BEA3BE93BE83BE73BE63BE53BE4",
		x"FFFFFFFFFFFFFFFF3BFF3BFE3BFD3BFC3BFB3BFA3BF93BF83BF73BF63BF53BF4",
		x"3C0F3C0E3C0D3C0C3C0B3C0A3C093C083C073C063C053C043C033C023C013C00",
		x"3C1F3C1E3C1D3C1C3C1B3C1A3C193C183C173C163C153C143C133C123C113C10",
		x"3C2F3C2E3C2D3C2C3C2B3C2A3C293C283C273C263C253C243C233C223C213C20",
		x"3C3F3C3E3C3D3C3C3C3B3C3A3C393C383C373C363C353C343C333C323C313C30",
		x"3C4B3C4A3C493C483C473C463C453C443C433C423C413C40FFFFFFFFFFFFFFFF",
		x"3C5B3C5A3C593C583C573C563C553C543C533C523C513C503C4F3C4E3C4D3C4C",
		x"3C6B3C6A3C693C683C673C663C653C643C633C623C613C603C5F3C5E3C5D3C5C",
		x"3C7B3C7A3C793C783C773C763C753C743C733C723C713C703C6F3C6E3C6D3C6C",
		x"3C873C863C853C843C833C823C813C80FFFFFFFFFFFFFFFF3C7F3C7E3C7D3C7C",
		x"3C973C963C953C943C933C923C913C903C8F3C8E3C8D3C8C3C8B3C8A3C893C88",
		x"3CA73CA63CA53CA43CA33CA23CA13CA03C9F3C9E3C9D3C9C3C9B3C9A3C993C98",
		x"3CB73CB63CB53CB43CB33CB23CB13CB03CAF3CAE3CAD3CAC3CAB3CAA3CA93CA8",
		x"3CC33CC23CC13CC0FFFFFFFFFFFFFFFF3CBF3CBE3CBD3CBC3CBB3CBA3CB93CB8",
		x"3CD33CD23CD13CD03CCF3CCE3CCD3CCC3CCB3CCA3CC93CC83CC73CC63CC53CC4",
		x"3CE33CE23CE13CE03CDF3CDE3CDD3CDC3CDB3CDA3CD93CD83CD73CD63CD53CD4",
		x"3CF33CF23CF13CF03CEF3CEE3CED3CEC3CEB3CEA3CE93CE83CE73CE63CE53CE4",
		x"FFFFFFFFFFFFFFFF3CFF3CFE3CFD3CFC3CFB3CFA3CF93CF83CF73CF63CF53CF4",
		x"3D0F3D0E3D0D3D0C3D0B3D0A3D093D083D073D063D053D043D033D023D013D00",
		x"3D1F3D1E3D1D3D1C3D1B3D1A3D193D183D173D163D153D143D133D123D113D10",
		x"3D2F3D2E3D2D3D2C3D2B3D2A3D293D283D273D263D253D243D233D223D213D20",
		x"3D3F3D3E3D3D3D3C3D3B3D3A3D393D383D373D363D353D343D333D323D313D30",
		x"3D4B3D4A3D493D483D473D463D453D443D433D423D413D40FFFFFFFFFFFFFFFF",
		x"3D5B3D5A3D593D583D573D563D553D543D533D523D513D503D4F3D4E3D4D3D4C",
		x"3D6B3D6A3D693D683D673D663D653D643D633D623D613D603D5F3D5E3D5D3D5C",
		x"3D7B3D7A3D793D783D773D763D753D743D733D723D713D703D6F3D6E3D6D3D6C",
		x"3D873D863D853D843D833D823D813D80FFFFFFFFFFFFFFFF3D7F3D7E3D7D3D7C",
		x"3D973D963D953D943D933D923D913D903D8F3D8E3D8D3D8C3D8B3D8A3D893D88",
		x"3DA73DA63DA53DA43DA33DA23DA13DA03D9F3D9E3D9D3D9C3D9B3D9A3D993D98",
		x"3DB73DB63DB53DB43DB33DB23DB13DB03DAF3DAE3DAD3DAC3DAB3DAA3DA93DA8",
		x"3DC33DC23DC13DC0FFFFFFFFFFFFFFFF3DBF3DBE3DBD3DBC3DBB3DBA3DB93DB8",
		x"3DD33DD23DD13DD03DCF3DCE3DCD3DCC3DCB3DCA3DC93DC83DC73DC63DC53DC4",
		x"3DE33DE23DE13DE03DDF3DDE3DDD3DDC3DDB3DDA3DD93DD83DD73DD63DD53DD4",
		x"3DF33DF23DF13DF03DEF3DEE3DED3DEC3DEB3DEA3DE93DE83DE73DE63DE53DE4",
		x"FFFFFFFFFFFFFFFF3DFF3DFE3DFD3DFC3DFB3DFA3DF93DF83DF73DF63DF53DF4",
		x"3E0F3E0E3E0D3E0C3E0B3E0A3E093E083E073E063E053E043E033E023E013E00",
		x"3E1F3E1E3E1D3E1C3E1B3E1A3E193E183E173E163E153E143E133E123E113E10",
		x"3E2F3E2E3E2D3E2C3E2B3E2A3E293E283E273E263E253E243E233E223E213E20",
		x"3E3F3E3E3E3D3E3C3E3B3E3A3E393E383E373E363E353E343E333E323E313E30",
		x"3E4B3E4A3E493E483E473E463E453E443E433E423E413E40FFFFFFFFFFFFFFFF",
		x"3E5B3E5A3E593E583E573E563E553E543E533E523E513E503E4F3E4E3E4D3E4C",
		x"3E6B3E6A3E693E683E673E663E653E643E633E623E613E603E5F3E5E3E5D3E5C",
		x"3E7B3E7A3E793E783E773E763E753E743E733E723E713E703E6F3E6E3E6D3E6C",
		x"3E873E863E853E843E833E823E813E80FFFFFFFFFFFFFFFF3E7F3E7E3E7D3E7C",
		x"3E973E963E953E943E933E923E913E903E8F3E8E3E8D3E8C3E8B3E8A3E893E88",
		x"3EA73EA63EA53EA43EA33EA23EA13EA03E9F3E9E3E9D3E9C3E9B3E9A3E993E98",
		x"3EB73EB63EB53EB43EB33EB23EB13EB03EAF3EAE3EAD3EAC3EAB3EAA3EA93EA8",
		x"3EC33EC23EC13EC0FFFFFFFFFFFFFFFF3EBF3EBE3EBD3EBC3EBB3EBA3EB93EB8",
		x"3ED33ED23ED13ED03ECF3ECE3ECD3ECC3ECB3ECA3EC93EC83EC73EC63EC53EC4",
		x"3EE33EE23EE13EE03EDF3EDE3EDD3EDC3EDB3EDA3ED93ED83ED73ED63ED53ED4",
		x"3EF33EF23EF13EF03EEF3EEE3EED3EEC3EEB3EEA3EE93EE83EE73EE63EE53EE4",
		x"FFFFFFFFFFFFFFFF3EFF3EFE3EFD3EFC3EFB3EFA3EF93EF83EF73EF63EF53EF4",
		x"3F0F3F0E3F0D3F0C3F0B3F0A3F093F083F073F063F053F043F033F023F013F00",
		x"3F1F3F1E3F1D3F1C3F1B3F1A3F193F183F173F163F153F143F133F123F113F10",
		x"3F2F3F2E3F2D3F2C3F2B3F2A3F293F283F273F263F253F243F233F223F213F20",
		x"3F3F3F3E3F3D3F3C3F3B3F3A3F393F383F373F363F353F343F333F323F313F30",
		x"3F4B3F4A3F493F483F473F463F453F443F433F423F413F40FFFFFFFFFFFFFFFF",
		x"3F5B3F5A3F593F583F573F563F553F543F533F523F513F503F4F3F4E3F4D3F4C",
		x"3F6B3F6A3F693F683F673F663F653F643F633F623F613F603F5F3F5E3F5D3F5C",
		x"3F7B3F7A3F793F783F773F763F753F743F733F723F713F703F6F3F6E3F6D3F6C",
		x"3F873F863F853F843F833F823F813F80FFFFFFFFFFFFFFFF3F7F3F7E3F7D3F7C",
		x"3F973F963F953F943F933F923F913F903F8F3F8E3F8D3F8C3F8B3F8A3F893F88",
		x"3FA73FA63FA53FA43FA33FA23FA13FA03F9F3F9E3F9D3F9C3F9B3F9A3F993F98",
		x"3FB73FB63FB53FB43FB33FB23FB13FB03FAF3FAE3FAD3FAC3FAB3FAA3FA93FA8",
		x"3FC33FC23FC13FC0FFFFFFFFFFFFFFFF3FBF3FBE3FBD3FBC3FBB3FBA3FB93FB8",
		x"3FD33FD23FD13FD03FCF3FCE3FCD3FCC3FCB3FCA3FC93FC83FC73FC63FC53FC4",
		x"3FE33FE23FE13FE03FDF3FDE3FDD3FDC3FDB3FDA3FD93FD83FD73FD63FD53FD4",
		x"3FF33FF23FF13FF03FEF3FEE3FED3FEC3FEB3FEA3FE93FE83FE73FE63FE53FE4",
		x"FFFFFFFFFFFFFFFF3FFF3FFE3FFD3FFC3FFB3FFA3FF93FF83FF73FF63FF53FF4",
		x"400F400E400D400C400B400A4009400840074006400540044003400240014000",
		x"401F401E401D401C401B401A4019401840174016401540144013401240114010",
		x"402F402E402D402C402B402A4029402840274026402540244023402240214020",
		x"403F403E403D403C403B403A4039403840374036403540344033403240314030",
		x"404B404A4049404840474046404540444043404240414040FFFFFFFFFFFFFFFF",
		x"405B405A4059405840574056405540544053405240514050404F404E404D404C",
		x"406B406A4069406840674066406540644063406240614060405F405E405D405C",
		x"407B407A4079407840774076407540744073407240714070406F406E406D406C",
		x"40874086408540844083408240814080FFFFFFFFFFFFFFFF407F407E407D407C",
		x"40974096409540944093409240914090408F408E408D408C408B408A40894088",
		x"40A740A640A540A440A340A240A140A0409F409E409D409C409B409A40994098",
		x"40B740B640B540B440B340B240B140B040AF40AE40AD40AC40AB40AA40A940A8",
		x"40C340C240C140C0FFFFFFFFFFFFFFFF40BF40BE40BD40BC40BB40BA40B940B8",
		x"40D340D240D140D040CF40CE40CD40CC40CB40CA40C940C840C740C640C540C4",
		x"40E340E240E140E040DF40DE40DD40DC40DB40DA40D940D840D740D640D540D4",
		x"40F340F240F140F040EF40EE40ED40EC40EB40EA40E940E840E740E640E540E4",
		x"FFFFFFFFFFFFFFFF40FF40FE40FD40FC40FB40FA40F940F840F740F640F540F4",
		x"410F410E410D410C410B410A4109410841074106410541044103410241014100",
		x"411F411E411D411C411B411A4119411841174116411541144113411241114110",
		x"412F412E412D412C412B412A4129412841274126412541244123412241214120",
		x"413F413E413D413C413B413A4139413841374136413541344133413241314130",
		x"414B414A4149414841474146414541444143414241414140FFFFFFFFFFFFFFFF",
		x"415B415A4159415841574156415541544153415241514150414F414E414D414C",
		x"416B416A4169416841674166416541644163416241614160415F415E415D415C",
		x"417B417A4179417841774176417541744173417241714170416F416E416D416C",
		x"41874186418541844183418241814180FFFFFFFFFFFFFFFF417F417E417D417C",
		x"41974196419541944193419241914190418F418E418D418C418B418A41894188",
		x"41A741A641A541A441A341A241A141A0419F419E419D419C419B419A41994198",
		x"41B741B641B541B441B341B241B141B041AF41AE41AD41AC41AB41AA41A941A8",
		x"41C341C241C141C0FFFFFFFFFFFFFFFF41BF41BE41BD41BC41BB41BA41B941B8",
		x"41D341D241D141D041CF41CE41CD41CC41CB41CA41C941C841C741C641C541C4",
		x"41E341E241E141E041DF41DE41DD41DC41DB41DA41D941D841D741D641D541D4",
		x"41F341F241F141F041EF41EE41ED41EC41EB41EA41E941E841E741E641E541E4",
		x"FFFFFFFFFFFFFFFF41FF41FE41FD41FC41FB41FA41F941F841F741F641F541F4",
		x"420F420E420D420C420B420A4209420842074206420542044203420242014200",
		x"421F421E421D421C421B421A4219421842174216421542144213421242114210",
		x"422F422E422D422C422B422A4229422842274226422542244223422242214220",
		x"423F423E423D423C423B423A4239423842374236423542344233423242314230",
		x"424B424A4249424842474246424542444243424242414240FFFFFFFFFFFFFFFF",
		x"425B425A4259425842574256425542544253425242514250424F424E424D424C",
		x"426B426A4269426842674266426542644263426242614260425F425E425D425C",
		x"427B427A4279427842774276427542744273427242714270426F426E426D426C",
		x"42874286428542844283428242814280FFFFFFFFFFFFFFFF427F427E427D427C",
		x"42974296429542944293429242914290428F428E428D428C428B428A42894288",
		x"42A742A642A542A442A342A242A142A0429F429E429D429C429B429A42994298",
		x"42B742B642B542B442B342B242B142B042AF42AE42AD42AC42AB42AA42A942A8",
		x"42C342C242C142C0FFFFFFFFFFFFFFFF42BF42BE42BD42BC42BB42BA42B942B8",
		x"42D342D242D142D042CF42CE42CD42CC42CB42CA42C942C842C742C642C542C4",
		x"42E342E242E142E042DF42DE42DD42DC42DB42DA42D942D842D742D642D542D4",
		x"42F342F242F142F042EF42EE42ED42EC42EB42EA42E942E842E742E642E542E4",
		x"FFFFFFFFFFFFFFFF42FF42FE42FD42FC42FB42FA42F942F842F742F642F542F4",
		x"430F430E430D430C430B430A4309430843074306430543044303430243014300",
		x"431F431E431D431C431B431A4319431843174316431543144313431243114310",
		x"432F432E432D432C432B432A4329432843274326432543244323432243214320",
		x"433F433E433D433C433B433A4339433843374336433543344333433243314330",
		x"434B434A4349434843474346434543444343434243414340FFFFFFFFFFFFFFFF",
		x"435B435A4359435843574356435543544353435243514350434F434E434D434C",
		x"436B436A4369436843674366436543644363436243614360435F435E435D435C",
		x"437B437A4379437843774376437543744373437243714370436F436E436D436C",
		x"43874386438543844383438243814380FFFFFFFFFFFFFFFF437F437E437D437C",
		x"43974396439543944393439243914390438F438E438D438C438B438A43894388",
		x"43A743A643A543A443A343A243A143A0439F439E439D439C439B439A43994398",
		x"43B743B643B543B443B343B243B143B043AF43AE43AD43AC43AB43AA43A943A8",
		x"43C343C243C143C0FFFFFFFFFFFFFFFF43BF43BE43BD43BC43BB43BA43B943B8",
		x"43D343D243D143D043CF43CE43CD43CC43CB43CA43C943C843C743C643C543C4",
		x"43E343E243E143E043DF43DE43DD43DC43DB43DA43D943D843D743D643D543D4",
		x"43F343F243F143F043EF43EE43ED43EC43EB43EA43E943E843E743E643E543E4",
		x"FFFFFFFFFFFFFFFF43FF43FE43FD43FC43FB43FA43F943F843F743F643F543F4",
		x"440F440E440D440C440B440A4409440844074406440544044403440244014400",
		x"441F441E441D441C441B441A4419441844174416441544144413441244114410",
		x"442F442E442D442C442B442A4429442844274426442544244423442244214420",
		x"443F443E443D443C443B443A4439443844374436443544344433443244314430",
		x"444B444A4449444844474446444544444443444244414440FFFFFFFFFFFFFFFF",
		x"445B445A4459445844574456445544544453445244514450444F444E444D444C",
		x"446B446A4469446844674466446544644463446244614460445F445E445D445C",
		x"447B447A4479447844774476447544744473447244714470446F446E446D446C",
		x"44874486448544844483448244814480FFFFFFFFFFFFFFFF447F447E447D447C",
		x"44974496449544944493449244914490448F448E448D448C448B448A44894488",
		x"44A744A644A544A444A344A244A144A0449F449E449D449C449B449A44994498",
		x"44B744B644B544B444B344B244B144B044AF44AE44AD44AC44AB44AA44A944A8",
		x"44C344C244C144C0FFFFFFFFFFFFFFFF44BF44BE44BD44BC44BB44BA44B944B8",
		x"44D344D244D144D044CF44CE44CD44CC44CB44CA44C944C844C744C644C544C4",
		x"44E344E244E144E044DF44DE44DD44DC44DB44DA44D944D844D744D644D544D4",
		x"44F344F244F144F044EF44EE44ED44EC44EB44EA44E944E844E744E644E544E4",
		x"FFFFFFFFFFFFFFFF44FF44FE44FD44FC44FB44FA44F944F844F744F644F544F4",
		x"450F450E450D450C450B450A4509450845074506450545044503450245014500",
		x"451F451E451D451C451B451A4519451845174516451545144513451245114510",
		x"452F452E452D452C452B452A4529452845274526452545244523452245214520",
		x"453F453E453D453C453B453A4539453845374536453545344533453245314530",
		x"454B454A4549454845474546454545444543454245414540FFFFFFFFFFFFFFFF",
		x"455B455A4559455845574556455545544553455245514550454F454E454D454C",
		x"456B456A4569456845674566456545644563456245614560455F455E455D455C",
		x"457B457A4579457845774576457545744573457245714570456F456E456D456C",
		x"45874586458545844583458245814580FFFFFFFFFFFFFFFF457F457E457D457C",
		x"45974596459545944593459245914590458F458E458D458C458B458A45894588",
		x"45A745A645A545A445A345A245A145A0459F459E459D459C459B459A45994598",
		x"45B745B645B545B445B345B245B145B045AF45AE45AD45AC45AB45AA45A945A8",
		x"45C345C245C145C0FFFFFFFFFFFFFFFF45BF45BE45BD45BC45BB45BA45B945B8",
		x"45D345D245D145D045CF45CE45CD45CC45CB45CA45C945C845C745C645C545C4",
		x"45E345E245E145E045DF45DE45DD45DC45DB45DA45D945D845D745D645D545D4",
		x"45F345F245F145F045EF45EE45ED45EC45EB45EA45E945E845E745E645E545E4",
		x"FFFFFFFFFFFFFFFF45FF45FE45FD45FC45FB45FA45F945F845F745F645F545F4",
		x"460F460E460D460C460B460A4609460846074606460546044603460246014600",
		x"461F461E461D461C461B461A4619461846174616461546144613461246114610",
		x"462F462E462D462C462B462A4629462846274626462546244623462246214620",
		x"463F463E463D463C463B463A4639463846374636463546344633463246314630",
		x"464B464A4649464846474646464546444643464246414640FFFFFFFFFFFFFFFF",
		x"465B465A4659465846574656465546544653465246514650464F464E464D464C",
		x"466B466A4669466846674666466546644663466246614660465F465E465D465C",
		x"467B467A4679467846774676467546744673467246714670466F466E466D466C",
		x"46874686468546844683468246814680FFFFFFFFFFFFFFFF467F467E467D467C",
		x"46974696469546944693469246914690468F468E468D468C468B468A46894688",
		x"46A746A646A546A446A346A246A146A0469F469E469D469C469B469A46994698",
		x"46B746B646B546B446B346B246B146B046AF46AE46AD46AC46AB46AA46A946A8",
		x"46C346C246C146C0FFFFFFFFFFFFFFFF46BF46BE46BD46BC46BB46BA46B946B8",
		x"46D346D246D146D046CF46CE46CD46CC46CB46CA46C946C846C746C646C546C4",
		x"46E346E246E146E046DF46DE46DD46DC46DB46DA46D946D846D746D646D546D4",
		x"46F346F246F146F046EF46EE46ED46EC46EB46EA46E946E846E746E646E546E4",
		x"FFFFFFFFFFFFFFFF46FF46FE46FD46FC46FB46FA46F946F846F746F646F546F4",
		x"470F470E470D470C470B470A4709470847074706470547044703470247014700",
		x"471F471E471D471C471B471A4719471847174716471547144713471247114710",
		x"472F472E472D472C472B472A4729472847274726472547244723472247214720",
		x"473F473E473D473C473B473A4739473847374736473547344733473247314730",
		x"474B474A4749474847474746474547444743474247414740FFFFFFFFFFFFFFFF",
		x"475B475A4759475847574756475547544753475247514750474F474E474D474C",
		x"476B476A4769476847674766476547644763476247614760475F475E475D475C",
		x"477B477A4779477847774776477547744773477247714770476F476E476D476C",
		x"47874786478547844783478247814780FFFFFFFFFFFFFFFF477F477E477D477C",
		x"47974796479547944793479247914790478F478E478D478C478B478A47894788",
		x"47A747A647A547A447A347A247A147A0479F479E479D479C479B479A47994798",
		x"47B747B647B547B447B347B247B147B047AF47AE47AD47AC47AB47AA47A947A8",
		x"47C347C247C147C0FFFFFFFFFFFFFFFF47BF47BE47BD47BC47BB47BA47B947B8",
		x"47D347D247D147D047CF47CE47CD47CC47CB47CA47C947C847C747C647C547C4",
		x"47E347E247E147E047DF47DE47DD47DC47DB47DA47D947D847D747D647D547D4",
		x"47F347F247F147F047EF47EE47ED47EC47EB47EA47E947E847E747E647E547E4",
		x"FFFFFFFFFFFFFFFF47FF47FE47FD47FC47FB47FA47F947F847F747F647F547F4",
		x"480F480E480D480C480B480A4809480848074806480548044803480248014800",
		x"481F481E481D481C481B481A4819481848174816481548144813481248114810",
		x"482F482E482D482C482B482A4829482848274826482548244823482248214820",
		x"483F483E483D483C483B483A4839483848374836483548344833483248314830",
		x"484B484A4849484848474846484548444843484248414840FFFFFFFFFFFFFFFF",
		x"485B485A4859485848574856485548544853485248514850484F484E484D484C",
		x"486B486A4869486848674866486548644863486248614860485F485E485D485C",
		x"487B487A4879487848774876487548744873487248714870486F486E486D486C",
		x"48874886488548844883488248814880FFFFFFFFFFFFFFFF487F487E487D487C",
		x"48974896489548944893489248914890488F488E488D488C488B488A48894888",
		x"48A748A648A548A448A348A248A148A0489F489E489D489C489B489A48994898",
		x"48B748B648B548B448B348B248B148B048AF48AE48AD48AC48AB48AA48A948A8",
		x"48C348C248C148C0FFFFFFFFFFFFFFFF48BF48BE48BD48BC48BB48BA48B948B8",
		x"48D348D248D148D048CF48CE48CD48CC48CB48CA48C948C848C748C648C548C4",
		x"48E348E248E148E048DF48DE48DD48DC48DB48DA48D948D848D748D648D548D4",
		x"48F348F248F148F048EF48EE48ED48EC48EB48EA48E948E848E748E648E548E4",
		x"FFFFFFFFFFFFFFFF48FF48FE48FD48FC48FB48FA48F948F848F748F648F548F4",
		x"490F490E490D490C490B490A4909490849074906490549044903490249014900",
		x"491F491E491D491C491B491A4919491849174916491549144913491249114910",
		x"492F492E492D492C492B492A4929492849274926492549244923492249214920",
		x"493F493E493D493C493B493A4939493849374936493549344933493249314930",
		x"494B494A4949494849474946494549444943494249414940FFFFFFFFFFFFFFFF",
		x"495B495A4959495849574956495549544953495249514950494F494E494D494C",
		x"496B496A4969496849674966496549644963496249614960495F495E495D495C",
		x"497B497A4979497849774976497549744973497249714970496F496E496D496C",
		x"49874986498549844983498249814980FFFFFFFFFFFFFFFF497F497E497D497C",
		x"49974996499549944993499249914990498F498E498D498C498B498A49894988",
		x"49A749A649A549A449A349A249A149A0499F499E499D499C499B499A49994998",
		x"49B749B649B549B449B349B249B149B049AF49AE49AD49AC49AB49AA49A949A8",
		x"49C349C249C149C0FFFFFFFFFFFFFFFF49BF49BE49BD49BC49BB49BA49B949B8",
		x"49D349D249D149D049CF49CE49CD49CC49CB49CA49C949C849C749C649C549C4",
		x"49E349E249E149E049DF49DE49DD49DC49DB49DA49D949D849D749D649D549D4",
		x"49F349F249F149F049EF49EE49ED49EC49EB49EA49E949E849E749E649E549E4",
		x"FFFFFFFFFFFFFFFF49FF49FE49FD49FC49FB49FA49F949F849F749F649F549F4",
		x"4A0F4A0E4A0D4A0C4A0B4A0A4A094A084A074A064A054A044A034A024A014A00",
		x"4A1F4A1E4A1D4A1C4A1B4A1A4A194A184A174A164A154A144A134A124A114A10",
		x"4A2F4A2E4A2D4A2C4A2B4A2A4A294A284A274A264A254A244A234A224A214A20",
		x"4A3F4A3E4A3D4A3C4A3B4A3A4A394A384A374A364A354A344A334A324A314A30",
		x"4A4B4A4A4A494A484A474A464A454A444A434A424A414A40FFFFFFFFFFFFFFFF",
		x"4A5B4A5A4A594A584A574A564A554A544A534A524A514A504A4F4A4E4A4D4A4C",
		x"4A6B4A6A4A694A684A674A664A654A644A634A624A614A604A5F4A5E4A5D4A5C",
		x"4A7B4A7A4A794A784A774A764A754A744A734A724A714A704A6F4A6E4A6D4A6C",
		x"4A874A864A854A844A834A824A814A80FFFFFFFFFFFFFFFF4A7F4A7E4A7D4A7C",
		x"4A974A964A954A944A934A924A914A904A8F4A8E4A8D4A8C4A8B4A8A4A894A88",
		x"4AA74AA64AA54AA44AA34AA24AA14AA04A9F4A9E4A9D4A9C4A9B4A9A4A994A98",
		x"4AB74AB64AB54AB44AB34AB24AB14AB04AAF4AAE4AAD4AAC4AAB4AAA4AA94AA8",
		x"4AC34AC24AC14AC0FFFFFFFFFFFFFFFF4ABF4ABE4ABD4ABC4ABB4ABA4AB94AB8",
		x"4AD34AD24AD14AD04ACF4ACE4ACD4ACC4ACB4ACA4AC94AC84AC74AC64AC54AC4",
		x"4AE34AE24AE14AE04ADF4ADE4ADD4ADC4ADB4ADA4AD94AD84AD74AD64AD54AD4",
		x"4AF34AF24AF14AF04AEF4AEE4AED4AEC4AEB4AEA4AE94AE84AE74AE64AE54AE4",
		x"FFFFFFFFFFFFFFFF4AFF4AFE4AFD4AFC4AFB4AFA4AF94AF84AF74AF64AF54AF4",
		x"4B0F4B0E4B0D4B0C4B0B4B0A4B094B084B074B064B054B044B034B024B014B00",
		x"4B1F4B1E4B1D4B1C4B1B4B1A4B194B184B174B164B154B144B134B124B114B10",
		x"4B2F4B2E4B2D4B2C4B2B4B2A4B294B284B274B264B254B244B234B224B214B20",
		x"4B3F4B3E4B3D4B3C4B3B4B3A4B394B384B374B364B354B344B334B324B314B30",
		x"4B4B4B4A4B494B484B474B464B454B444B434B424B414B40FFFFFFFFFFFFFFFF",
		x"4B5B4B5A4B594B584B574B564B554B544B534B524B514B504B4F4B4E4B4D4B4C",
		x"4B6B4B6A4B694B684B674B664B654B644B634B624B614B604B5F4B5E4B5D4B5C",
		x"4B7B4B7A4B794B784B774B764B754B744B734B724B714B704B6F4B6E4B6D4B6C",
		x"4B874B864B854B844B834B824B814B80FFFFFFFFFFFFFFFF4B7F4B7E4B7D4B7C",
		x"4B974B964B954B944B934B924B914B904B8F4B8E4B8D4B8C4B8B4B8A4B894B88",
		x"4BA74BA64BA54BA44BA34BA24BA14BA04B9F4B9E4B9D4B9C4B9B4B9A4B994B98",
		x"4BB74BB64BB54BB44BB34BB24BB14BB04BAF4BAE4BAD4BAC4BAB4BAA4BA94BA8",
		x"4BC34BC24BC14BC0FFFFFFFFFFFFFFFF4BBF4BBE4BBD4BBC4BBB4BBA4BB94BB8",
		x"4BD34BD24BD14BD04BCF4BCE4BCD4BCC4BCB4BCA4BC94BC84BC74BC64BC54BC4",
		x"4BE34BE24BE14BE04BDF4BDE4BDD4BDC4BDB4BDA4BD94BD84BD74BD64BD54BD4",
		x"4BF34BF24BF14BF04BEF4BEE4BED4BEC4BEB4BEA4BE94BE84BE74BE64BE54BE4",
		x"FFFFFFFFFFFFFFFF4BFF4BFE4BFD4BFC4BFB4BFA4BF94BF84BF74BF64BF54BF4",
		x"4C0F4C0E4C0D4C0C4C0B4C0A4C094C084C074C064C054C044C034C024C014C00",
		x"4C1F4C1E4C1D4C1C4C1B4C1A4C194C184C174C164C154C144C134C124C114C10",
		x"4C2F4C2E4C2D4C2C4C2B4C2A4C294C284C274C264C254C244C234C224C214C20",
		x"4C3F4C3E4C3D4C3C4C3B4C3A4C394C384C374C364C354C344C334C324C314C30",
		x"4C4B4C4A4C494C484C474C464C454C444C434C424C414C40FFFFFFFFFFFFFFFF",
		x"4C5B4C5A4C594C584C574C564C554C544C534C524C514C504C4F4C4E4C4D4C4C",
		x"4C6B4C6A4C694C684C674C664C654C644C634C624C614C604C5F4C5E4C5D4C5C",
		x"4C7B4C7A4C794C784C774C764C754C744C734C724C714C704C6F4C6E4C6D4C6C",
		x"4C874C864C854C844C834C824C814C80FFFFFFFFFFFFFFFF4C7F4C7E4C7D4C7C",
		x"4C974C964C954C944C934C924C914C904C8F4C8E4C8D4C8C4C8B4C8A4C894C88",
		x"4CA74CA64CA54CA44CA34CA24CA14CA04C9F4C9E4C9D4C9C4C9B4C9A4C994C98",
		x"4CB74CB64CB54CB44CB34CB24CB14CB04CAF4CAE4CAD4CAC4CAB4CAA4CA94CA8",
		x"4CC34CC24CC14CC0FFFFFFFFFFFFFFFF4CBF4CBE4CBD4CBC4CBB4CBA4CB94CB8",
		x"4CD34CD24CD14CD04CCF4CCE4CCD4CCC4CCB4CCA4CC94CC84CC74CC64CC54CC4",
		x"4CE34CE24CE14CE04CDF4CDE4CDD4CDC4CDB4CDA4CD94CD84CD74CD64CD54CD4",
		x"4CF34CF24CF14CF04CEF4CEE4CED4CEC4CEB4CEA4CE94CE84CE74CE64CE54CE4",
		x"FFFFFFFFFFFFFFFF4CFF4CFE4CFD4CFC4CFB4CFA4CF94CF84CF74CF64CF54CF4",
		x"4D0F4D0E4D0D4D0C4D0B4D0A4D094D084D074D064D054D044D034D024D014D00",
		x"4D1F4D1E4D1D4D1C4D1B4D1A4D194D184D174D164D154D144D134D124D114D10",
		x"4D2F4D2E4D2D4D2C4D2B4D2A4D294D284D274D264D254D244D234D224D214D20",
		x"4D3F4D3E4D3D4D3C4D3B4D3A4D394D384D374D364D354D344D334D324D314D30",
		x"4D4B4D4A4D494D484D474D464D454D444D434D424D414D40FFFFFFFFFFFFFFFF",
		x"4D5B4D5A4D594D584D574D564D554D544D534D524D514D504D4F4D4E4D4D4D4C",
		x"4D6B4D6A4D694D684D674D664D654D644D634D624D614D604D5F4D5E4D5D4D5C",
		x"4D7B4D7A4D794D784D774D764D754D744D734D724D714D704D6F4D6E4D6D4D6C",
		x"4D874D864D854D844D834D824D814D80FFFFFFFFFFFFFFFF4D7F4D7E4D7D4D7C",
		x"4D974D964D954D944D934D924D914D904D8F4D8E4D8D4D8C4D8B4D8A4D894D88",
		x"4DA74DA64DA54DA44DA34DA24DA14DA04D9F4D9E4D9D4D9C4D9B4D9A4D994D98",
		x"4DB74DB64DB54DB44DB34DB24DB14DB04DAF4DAE4DAD4DAC4DAB4DAA4DA94DA8",
		x"4DC34DC24DC14DC0FFFFFFFFFFFFFFFF4DBF4DBE4DBD4DBC4DBB4DBA4DB94DB8",
		x"4DD34DD24DD14DD04DCF4DCE4DCD4DCC4DCB4DCA4DC94DC84DC74DC64DC54DC4",
		x"4DE34DE24DE14DE04DDF4DDE4DDD4DDC4DDB4DDA4DD94DD84DD74DD64DD54DD4",
		x"4DF34DF24DF14DF04DEF4DEE4DED4DEC4DEB4DEA4DE94DE84DE74DE64DE54DE4",
		x"FFFFFFFFFFFFFFFF4DFF4DFE4DFD4DFC4DFB4DFA4DF94DF84DF74DF64DF54DF4",
		x"4E0F4E0E4E0D4E0C4E0B4E0A4E094E084E074E064E054E044E034E024E014E00",
		x"4E1F4E1E4E1D4E1C4E1B4E1A4E194E184E174E164E154E144E134E124E114E10",
		x"4E2F4E2E4E2D4E2C4E2B4E2A4E294E284E274E264E254E244E234E224E214E20",
		x"4E3F4E3E4E3D4E3C4E3B4E3A4E394E384E374E364E354E344E334E324E314E30",
		x"4E4B4E4A4E494E484E474E464E454E444E434E424E414E40FFFFFFFFFFFFFFFF",
		x"4E5B4E5A4E594E584E574E564E554E544E534E524E514E504E4F4E4E4E4D4E4C",
		x"4E6B4E6A4E694E684E674E664E654E644E634E624E614E604E5F4E5E4E5D4E5C",
		x"4E7B4E7A4E794E784E774E764E754E744E734E724E714E704E6F4E6E4E6D4E6C",
		x"4E874E864E854E844E834E824E814E80FFFFFFFFFFFFFFFF4E7F4E7E4E7D4E7C",
		x"4E974E964E954E944E934E924E914E904E8F4E8E4E8D4E8C4E8B4E8A4E894E88",
		x"4EA74EA64EA54EA44EA34EA24EA14EA04E9F4E9E4E9D4E9C4E9B4E9A4E994E98",
		x"4EB74EB64EB54EB44EB34EB24EB14EB04EAF4EAE4EAD4EAC4EAB4EAA4EA94EA8",
		x"4EC34EC24EC14EC0FFFFFFFFFFFFFFFF4EBF4EBE4EBD4EBC4EBB4EBA4EB94EB8",
		x"4ED34ED24ED14ED04ECF4ECE4ECD4ECC4ECB4ECA4EC94EC84EC74EC64EC54EC4",
		x"4EE34EE24EE14EE04EDF4EDE4EDD4EDC4EDB4EDA4ED94ED84ED74ED64ED54ED4",
		x"4EF34EF24EF14EF04EEF4EEE4EED4EEC4EEB4EEA4EE94EE84EE74EE64EE54EE4",
		x"FFFFFFFFFFFFFFFF4EFF4EFE4EFD4EFC4EFB4EFA4EF94EF84EF74EF64EF54EF4",
		x"4F0F4F0E4F0D4F0C4F0B4F0A4F094F084F074F064F054F044F034F024F014F00",
		x"4F1F4F1E4F1D4F1C4F1B4F1A4F194F184F174F164F154F144F134F124F114F10",
		x"4F2F4F2E4F2D4F2C4F2B4F2A4F294F284F274F264F254F244F234F224F214F20",
		x"4F3F4F3E4F3D4F3C4F3B4F3A4F394F384F374F364F354F344F334F324F314F30",
		x"4F4B4F4A4F494F484F474F464F454F444F434F424F414F40FFFFFFFFFFFFFFFF",
		x"4F5B4F5A4F594F584F574F564F554F544F534F524F514F504F4F4F4E4F4D4F4C",
		x"4F6B4F6A4F694F684F674F664F654F644F634F624F614F604F5F4F5E4F5D4F5C",
		x"4F7B4F7A4F794F784F774F764F754F744F734F724F714F704F6F4F6E4F6D4F6C",
		x"4F874F864F854F844F834F824F814F80FFFFFFFFFFFFFFFF4F7F4F7E4F7D4F7C",
		x"4F974F964F954F944F934F924F914F904F8F4F8E4F8D4F8C4F8B4F8A4F894F88",
		x"4FA74FA64FA54FA44FA34FA24FA14FA04F9F4F9E4F9D4F9C4F9B4F9A4F994F98",
		x"4FB74FB64FB54FB44FB34FB24FB14FB04FAF4FAE4FAD4FAC4FAB4FAA4FA94FA8",
		x"4FC34FC24FC14FC0FFFFFFFFFFFFFFFF4FBF4FBE4FBD4FBC4FBB4FBA4FB94FB8",
		x"4FD34FD24FD14FD04FCF4FCE4FCD4FCC4FCB4FCA4FC94FC84FC74FC64FC54FC4",
		x"4FE34FE24FE14FE04FDF4FDE4FDD4FDC4FDB4FDA4FD94FD84FD74FD64FD54FD4",
		x"4FF34FF24FF14FF04FEF4FEE4FED4FEC4FEB4FEA4FE94FE84FE74FE64FE54FE4",
		x"FFFFFFFFFFFFFFFF4FFF4FFE4FFD4FFC4FFB4FFA4FF94FF84FF74FF64FF54FF4",
		x"500F500E500D500C500B500A5009500850075006500550045003500250015000",
		x"501F501E501D501C501B501A5019501850175016501550145013501250115010",
		x"502F502E502D502C502B502A5029502850275026502550245023502250215020",
		x"503F503E503D503C503B503A5039503850375036503550345033503250315030",
		x"504B504A5049504850475046504550445043504250415040FFFFFFFFFFFFFFFF",
		x"505B505A5059505850575056505550545053505250515050504F504E504D504C",
		x"506B506A5069506850675066506550645063506250615060505F505E505D505C",
		x"507B507A5079507850775076507550745073507250715070506F506E506D506C",
		x"50875086508550845083508250815080FFFFFFFFFFFFFFFF507F507E507D507C",
		x"50975096509550945093509250915090508F508E508D508C508B508A50895088",
		x"50A750A650A550A450A350A250A150A0509F509E509D509C509B509A50995098",
		x"50B750B650B550B450B350B250B150B050AF50AE50AD50AC50AB50AA50A950A8",
		x"50C350C250C150C0FFFFFFFFFFFFFFFF50BF50BE50BD50BC50BB50BA50B950B8",
		x"50D350D250D150D050CF50CE50CD50CC50CB50CA50C950C850C750C650C550C4",
		x"50E350E250E150E050DF50DE50DD50DC50DB50DA50D950D850D750D650D550D4",
		x"50F350F250F150F050EF50EE50ED50EC50EB50EA50E950E850E750E650E550E4",
		x"FFFFFFFFFFFFFFFF50FF50FE50FD50FC50FB50FA50F950F850F750F650F550F4",
		x"510F510E510D510C510B510A5109510851075106510551045103510251015100",
		x"511F511E511D511C511B511A5119511851175116511551145113511251115110",
		x"512F512E512D512C512B512A5129512851275126512551245123512251215120",
		x"513F513E513D513C513B513A5139513851375136513551345133513251315130",
		x"514B514A5149514851475146514551445143514251415140FFFFFFFFFFFFFFFF",
		x"515B515A5159515851575156515551545153515251515150514F514E514D514C",
		x"516B516A5169516851675166516551645163516251615160515F515E515D515C",
		x"517B517A5179517851775176517551745173517251715170516F516E516D516C",
		x"51875186518551845183518251815180FFFFFFFFFFFFFFFF517F517E517D517C",
		x"51975196519551945193519251915190518F518E518D518C518B518A51895188",
		x"51A751A651A551A451A351A251A151A0519F519E519D519C519B519A51995198",
		x"51B751B651B551B451B351B251B151B051AF51AE51AD51AC51AB51AA51A951A8",
		x"51C351C251C151C0FFFFFFFFFFFFFFFF51BF51BE51BD51BC51BB51BA51B951B8",
		x"51D351D251D151D051CF51CE51CD51CC51CB51CA51C951C851C751C651C551C4",
		x"51E351E251E151E051DF51DE51DD51DC51DB51DA51D951D851D751D651D551D4",
		x"51F351F251F151F051EF51EE51ED51EC51EB51EA51E951E851E751E651E551E4",
		x"FFFFFFFFFFFFFFFF51FF51FE51FD51FC51FB51FA51F951F851F751F651F551F4",
		x"520F520E520D520C520B520A5209520852075206520552045203520252015200",
		x"521F521E521D521C521B521A5219521852175216521552145213521252115210",
		x"522F522E522D522C522B522A5229522852275226522552245223522252215220",
		x"523F523E523D523C523B523A5239523852375236523552345233523252315230",
		x"524B524A5249524852475246524552445243524252415240FFFFFFFFFFFFFFFF",
		x"525B525A5259525852575256525552545253525252515250524F524E524D524C",
		x"526B526A5269526852675266526552645263526252615260525F525E525D525C",
		x"527B527A5279527852775276527552745273527252715270526F526E526D526C",
		x"52875286528552845283528252815280FFFFFFFFFFFFFFFF527F527E527D527C",
		x"52975296529552945293529252915290528F528E528D528C528B528A52895288",
		x"52A752A652A552A452A352A252A152A0529F529E529D529C529B529A52995298",
		x"52B752B652B552B452B352B252B152B052AF52AE52AD52AC52AB52AA52A952A8",
		x"52C352C252C152C0FFFFFFFFFFFFFFFF52BF52BE52BD52BC52BB52BA52B952B8",
		x"52D352D252D152D052CF52CE52CD52CC52CB52CA52C952C852C752C652C552C4",
		x"52E352E252E152E052DF52DE52DD52DC52DB52DA52D952D852D752D652D552D4",
		x"52F352F252F152F052EF52EE52ED52EC52EB52EA52E952E852E752E652E552E4",
		x"FFFFFFFFFFFFFFFF52FF52FE52FD52FC52FB52FA52F952F852F752F652F552F4",
		x"530F530E530D530C530B530A5309530853075306530553045303530253015300",
		x"531F531E531D531C531B531A5319531853175316531553145313531253115310",
		x"532F532E532D532C532B532A5329532853275326532553245323532253215320",
		x"533F533E533D533C533B533A5339533853375336533553345333533253315330",
		x"534B534A5349534853475346534553445343534253415340FFFFFFFFFFFFFFFF",
		x"535B535A5359535853575356535553545353535253515350534F534E534D534C",
		x"536B536A5369536853675366536553645363536253615360535F535E535D535C",
		x"537B537A5379537853775376537553745373537253715370536F536E536D536C",
		x"53875386538553845383538253815380FFFFFFFFFFFFFFFF537F537E537D537C",
		x"53975396539553945393539253915390538F538E538D538C538B538A53895388",
		x"53A753A653A553A453A353A253A153A0539F539E539D539C539B539A53995398",
		x"53B753B653B553B453B353B253B153B053AF53AE53AD53AC53AB53AA53A953A8",
		x"53C353C253C153C0FFFFFFFFFFFFFFFF53BF53BE53BD53BC53BB53BA53B953B8",
		x"53D353D253D153D053CF53CE53CD53CC53CB53CA53C953C853C753C653C553C4",
		x"53E353E253E153E053DF53DE53DD53DC53DB53DA53D953D853D753D653D553D4",
		x"53F353F253F153F053EF53EE53ED53EC53EB53EA53E953E853E753E653E553E4",
		x"FFFFFFFFFFFFFFFF53FF53FE53FD53FC53FB53FA53F953F853F753F653F553F4",
		x"540F540E540D540C540B540A5409540854075406540554045403540254015400",
		x"541F541E541D541C541B541A5419541854175416541554145413541254115410",
		x"542F542E542D542C542B542A5429542854275426542554245423542254215420",
		x"543F543E543D543C543B543A5439543854375436543554345433543254315430",
		x"544B544A5449544854475446544554445443544254415440FFFFFFFFFFFFFFFF",
		x"545B545A5459545854575456545554545453545254515450544F544E544D544C",
		x"546B546A5469546854675466546554645463546254615460545F545E545D545C",
		x"547B547A5479547854775476547554745473547254715470546F546E546D546C",
		x"54875486548554845483548254815480FFFFFFFFFFFFFFFF547F547E547D547C",
		x"54975496549554945493549254915490548F548E548D548C548B548A54895488",
		x"54A754A654A554A454A354A254A154A0549F549E549D549C549B549A54995498",
		x"54B754B654B554B454B354B254B154B054AF54AE54AD54AC54AB54AA54A954A8",
		x"54C354C254C154C0FFFFFFFFFFFFFFFF54BF54BE54BD54BC54BB54BA54B954B8",
		x"54D354D254D154D054CF54CE54CD54CC54CB54CA54C954C854C754C654C554C4",
		x"54E354E254E154E054DF54DE54DD54DC54DB54DA54D954D854D754D654D554D4",
		x"54F354F254F154F054EF54EE54ED54EC54EB54EA54E954E854E754E654E554E4",
		x"FFFFFFFFFFFFFFFF54FF54FE54FD54FC54FB54FA54F954F854F754F654F554F4",
		x"550F550E550D550C550B550A5509550855075506550555045503550255015500",
		x"551F551E551D551C551B551A5519551855175516551555145513551255115510",
		x"552F552E552D552C552B552A5529552855275526552555245523552255215520",
		x"553F553E553D553C553B553A5539553855375536553555345533553255315530",
		x"554B554A5549554855475546554555445543554255415540FFFFFFFFFFFFFFFF",
		x"555B555A5559555855575556555555545553555255515550554F554E554D554C",
		x"556B556A5569556855675566556555645563556255615560555F555E555D555C",
		x"557B557A5579557855775576557555745573557255715570556F556E556D556C",
		x"55875586558555845583558255815580FFFFFFFFFFFFFFFF557F557E557D557C",
		x"55975596559555945593559255915590558F558E558D558C558B558A55895588",
		x"55A755A655A555A455A355A255A155A0559F559E559D559C559B559A55995598",
		x"55B755B655B555B455B355B255B155B055AF55AE55AD55AC55AB55AA55A955A8",
		x"55C355C255C155C0FFFFFFFFFFFFFFFF55BF55BE55BD55BC55BB55BA55B955B8",
		x"55D355D255D155D055CF55CE55CD55CC55CB55CA55C955C855C755C655C555C4",
		x"55E355E255E155E055DF55DE55DD55DC55DB55DA55D955D855D755D655D555D4",
		x"55F355F255F155F055EF55EE55ED55EC55EB55EA55E955E855E755E655E555E4",
		x"FFFFFFFFFFFFFFFF55FF55FE55FD55FC55FB55FA55F955F855F755F655F555F4",
		x"560F560E560D560C560B560A5609560856075606560556045603560256015600",
		x"561F561E561D561C561B561A5619561856175616561556145613561256115610",
		x"562F562E562D562C562B562A5629562856275626562556245623562256215620",
		x"563F563E563D563C563B563A5639563856375636563556345633563256315630",
		x"564B564A5649564856475646564556445643564256415640FFFFFFFFFFFFFFFF",
		x"565B565A5659565856575656565556545653565256515650564F564E564D564C",
		x"566B566A5669566856675666566556645663566256615660565F565E565D565C",
		x"567B567A5679567856775676567556745673567256715670566F566E566D566C",
		x"56875686568556845683568256815680FFFFFFFFFFFFFFFF567F567E567D567C",
		x"56975696569556945693569256915690568F568E568D568C568B568A56895688",
		x"56A756A656A556A456A356A256A156A0569F569E569D569C569B569A56995698",
		x"56B756B656B556B456B356B256B156B056AF56AE56AD56AC56AB56AA56A956A8",
		x"56C356C256C156C0FFFFFFFFFFFFFFFF56BF56BE56BD56BC56BB56BA56B956B8",
		x"56D356D256D156D056CF56CE56CD56CC56CB56CA56C956C856C756C656C556C4",
		x"56E356E256E156E056DF56DE56DD56DC56DB56DA56D956D856D756D656D556D4",
		x"56F356F256F156F056EF56EE56ED56EC56EB56EA56E956E856E756E656E556E4",
		x"FFFFFFFFFFFFFFFF56FF56FE56FD56FC56FB56FA56F956F856F756F656F556F4",
		x"570F570E570D570C570B570A5709570857075706570557045703570257015700",
		x"571F571E571D571C571B571A5719571857175716571557145713571257115710",
		x"572F572E572D572C572B572A5729572857275726572557245723572257215720",
		x"573F573E573D573C573B573A5739573857375736573557345733573257315730",
		x"574B574A5749574857475746574557445743574257415740FFFFFFFFFFFFFFFF",
		x"575B575A5759575857575756575557545753575257515750574F574E574D574C",
		x"576B576A5769576857675766576557645763576257615760575F575E575D575C",
		x"577B577A5779577857775776577557745773577257715770576F576E576D576C",
		x"57875786578557845783578257815780FFFFFFFFFFFFFFFF577F577E577D577C",
		x"57975796579557945793579257915790578F578E578D578C578B578A57895788",
		x"57A757A657A557A457A357A257A157A0579F579E579D579C579B579A57995798",
		x"57B757B657B557B457B357B257B157B057AF57AE57AD57AC57AB57AA57A957A8",
		x"57C357C257C157C0FFFFFFFFFFFFFFFF57BF57BE57BD57BC57BB57BA57B957B8",
		x"57D357D257D157D057CF57CE57CD57CC57CB57CA57C957C857C757C657C557C4",
		x"57E357E257E157E057DF57DE57DD57DC57DB57DA57D957D857D757D657D557D4",
		x"57F357F257F157F057EF57EE57ED57EC57EB57EA57E957E857E757E657E557E4",
		x"FFFFFFFFFFFFFFFF57FF57FE57FD57FC57FB57FA57F957F857F757F657F557F4",
		x"580F580E580D580C580B580A5809580858075806580558045803580258015800",
		x"581F581E581D581C581B581A5819581858175816581558145813581258115810",
		x"582F582E582D582C582B582A5829582858275826582558245823582258215820",
		x"583F583E583D583C583B583A5839583858375836583558345833583258315830",
		x"584B584A5849584858475846584558445843584258415840FFFFFFFFFFFFFFFF",
		x"585B585A5859585858575856585558545853585258515850584F584E584D584C",
		x"586B586A5869586858675866586558645863586258615860585F585E585D585C",
		x"587B587A5879587858775876587558745873587258715870586F586E586D586C",
		x"58875886588558845883588258815880FFFFFFFFFFFFFFFF587F587E587D587C",
		x"58975896589558945893589258915890588F588E588D588C588B588A58895888",
		x"58A758A658A558A458A358A258A158A0589F589E589D589C589B589A58995898",
		x"58B758B658B558B458B358B258B158B058AF58AE58AD58AC58AB58AA58A958A8",
		x"58C358C258C158C0FFFFFFFFFFFFFFFF58BF58BE58BD58BC58BB58BA58B958B8",
		x"58D358D258D158D058CF58CE58CD58CC58CB58CA58C958C858C758C658C558C4",
		x"58E358E258E158E058DF58DE58DD58DC58DB58DA58D958D858D758D658D558D4",
		x"58F358F258F158F058EF58EE58ED58EC58EB58EA58E958E858E758E658E558E4",
		x"FFFFFFFFFFFFFFFF58FF58FE58FD58FC58FB58FA58F958F858F758F658F558F4",
		x"590F590E590D590C590B590A5909590859075906590559045903590259015900",
		x"591F591E591D591C591B591A5919591859175916591559145913591259115910",
		x"592F592E592D592C592B592A5929592859275926592559245923592259215920",
		x"593F593E593D593C593B593A5939593859375936593559345933593259315930",
		x"594B594A5949594859475946594559445943594259415940FFFFFFFFFFFFFFFF",
		x"595B595A5959595859575956595559545953595259515950594F594E594D594C",
		x"596B596A5969596859675966596559645963596259615960595F595E595D595C",
		x"597B597A5979597859775976597559745973597259715970596F596E596D596C",
		x"59875986598559845983598259815980FFFFFFFFFFFFFFFF597F597E597D597C",
		x"59975996599559945993599259915990598F598E598D598C598B598A59895988",
		x"59A759A659A559A459A359A259A159A0599F599E599D599C599B599A59995998",
		x"59B759B659B559B459B359B259B159B059AF59AE59AD59AC59AB59AA59A959A8",
		x"59C359C259C159C0FFFFFFFFFFFFFFFF59BF59BE59BD59BC59BB59BA59B959B8",
		x"59D359D259D159D059CF59CE59CD59CC59CB59CA59C959C859C759C659C559C4",
		x"59E359E259E159E059DF59DE59DD59DC59DB59DA59D959D859D759D659D559D4",
		x"59F359F259F159F059EF59EE59ED59EC59EB59EA59E959E859E759E659E559E4",
		x"FFFFFFFFFFFFFFFF59FF59FE59FD59FC59FB59FA59F959F859F759F659F559F4",
		x"5A0F5A0E5A0D5A0C5A0B5A0A5A095A085A075A065A055A045A035A025A015A00",
		x"5A1F5A1E5A1D5A1C5A1B5A1A5A195A185A175A165A155A145A135A125A115A10",
		x"5A2F5A2E5A2D5A2C5A2B5A2A5A295A285A275A265A255A245A235A225A215A20",
		x"5A3F5A3E5A3D5A3C5A3B5A3A5A395A385A375A365A355A345A335A325A315A30",
		x"5A4B5A4A5A495A485A475A465A455A445A435A425A415A40FFFFFFFFFFFFFFFF",
		x"5A5B5A5A5A595A585A575A565A555A545A535A525A515A505A4F5A4E5A4D5A4C",
		x"5A6B5A6A5A695A685A675A665A655A645A635A625A615A605A5F5A5E5A5D5A5C",
		x"5A7B5A7A5A795A785A775A765A755A745A735A725A715A705A6F5A6E5A6D5A6C",
		x"5A875A865A855A845A835A825A815A80FFFFFFFFFFFFFFFF5A7F5A7E5A7D5A7C",
		x"5A975A965A955A945A935A925A915A905A8F5A8E5A8D5A8C5A8B5A8A5A895A88",
		x"5AA75AA65AA55AA45AA35AA25AA15AA05A9F5A9E5A9D5A9C5A9B5A9A5A995A98",
		x"5AB75AB65AB55AB45AB35AB25AB15AB05AAF5AAE5AAD5AAC5AAB5AAA5AA95AA8",
		x"5AC35AC25AC15AC0FFFFFFFFFFFFFFFF5ABF5ABE5ABD5ABC5ABB5ABA5AB95AB8",
		x"5AD35AD25AD15AD05ACF5ACE5ACD5ACC5ACB5ACA5AC95AC85AC75AC65AC55AC4",
		x"5AE35AE25AE15AE05ADF5ADE5ADD5ADC5ADB5ADA5AD95AD85AD75AD65AD55AD4",
		x"5AF35AF25AF15AF05AEF5AEE5AED5AEC5AEB5AEA5AE95AE85AE75AE65AE55AE4",
		x"FFFFFFFFFFFFFFFF5AFF5AFE5AFD5AFC5AFB5AFA5AF95AF85AF75AF65AF55AF4",
		x"5B0F5B0E5B0D5B0C5B0B5B0A5B095B085B075B065B055B045B035B025B015B00",
		x"5B1F5B1E5B1D5B1C5B1B5B1A5B195B185B175B165B155B145B135B125B115B10",
		x"5B2F5B2E5B2D5B2C5B2B5B2A5B295B285B275B265B255B245B235B225B215B20",
		x"5B3F5B3E5B3D5B3C5B3B5B3A5B395B385B375B365B355B345B335B325B315B30",
		x"5B4B5B4A5B495B485B475B465B455B445B435B425B415B40FFFFFFFFFFFFFFFF",
		x"5B5B5B5A5B595B585B575B565B555B545B535B525B515B505B4F5B4E5B4D5B4C",
		x"5B6B5B6A5B695B685B675B665B655B645B635B625B615B605B5F5B5E5B5D5B5C",
		x"5B7B5B7A5B795B785B775B765B755B745B735B725B715B705B6F5B6E5B6D5B6C",
		x"5B875B865B855B845B835B825B815B80FFFFFFFFFFFFFFFF5B7F5B7E5B7D5B7C",
		x"5B975B965B955B945B935B925B915B905B8F5B8E5B8D5B8C5B8B5B8A5B895B88",
		x"5BA75BA65BA55BA45BA35BA25BA15BA05B9F5B9E5B9D5B9C5B9B5B9A5B995B98",
		x"5BB75BB65BB55BB45BB35BB25BB15BB05BAF5BAE5BAD5BAC5BAB5BAA5BA95BA8",
		x"5BC35BC25BC15BC0FFFFFFFFFFFFFFFF5BBF5BBE5BBD5BBC5BBB5BBA5BB95BB8",
		x"5BD35BD25BD15BD05BCF5BCE5BCD5BCC5BCB5BCA5BC95BC85BC75BC65BC55BC4",
		x"5BE35BE25BE15BE05BDF5BDE5BDD5BDC5BDB5BDA5BD95BD85BD75BD65BD55BD4",
		x"5BF35BF25BF15BF05BEF5BEE5BED5BEC5BEB5BEA5BE95BE85BE75BE65BE55BE4",
		x"FFFFFFFFFFFFFFFF5BFF5BFE5BFD5BFC5BFB5BFA5BF95BF85BF75BF65BF55BF4",
		x"5C0F5C0E5C0D5C0C5C0B5C0A5C095C085C075C065C055C045C035C025C015C00",
		x"5C1F5C1E5C1D5C1C5C1B5C1A5C195C185C175C165C155C145C135C125C115C10",
		x"5C2F5C2E5C2D5C2C5C2B5C2A5C295C285C275C265C255C245C235C225C215C20",
		x"5C3F5C3E5C3D5C3C5C3B5C3A5C395C385C375C365C355C345C335C325C315C30",
		x"5C4B5C4A5C495C485C475C465C455C445C435C425C415C40FFFFFFFFFFFFFFFF",
		x"5C5B5C5A5C595C585C575C565C555C545C535C525C515C505C4F5C4E5C4D5C4C",
		x"5C6B5C6A5C695C685C675C665C655C645C635C625C615C605C5F5C5E5C5D5C5C",
		x"5C7B5C7A5C795C785C775C765C755C745C735C725C715C705C6F5C6E5C6D5C6C",
		x"5C875C865C855C845C835C825C815C80FFFFFFFFFFFFFFFF5C7F5C7E5C7D5C7C",
		x"5C975C965C955C945C935C925C915C905C8F5C8E5C8D5C8C5C8B5C8A5C895C88",
		x"5CA75CA65CA55CA45CA35CA25CA15CA05C9F5C9E5C9D5C9C5C9B5C9A5C995C98",
		x"5CB75CB65CB55CB45CB35CB25CB15CB05CAF5CAE5CAD5CAC5CAB5CAA5CA95CA8",
		x"5CC35CC25CC15CC0FFFFFFFFFFFFFFFF5CBF5CBE5CBD5CBC5CBB5CBA5CB95CB8",
		x"5CD35CD25CD15CD05CCF5CCE5CCD5CCC5CCB5CCA5CC95CC85CC75CC65CC55CC4",
		x"5CE35CE25CE15CE05CDF5CDE5CDD5CDC5CDB5CDA5CD95CD85CD75CD65CD55CD4",
		x"5CF35CF25CF15CF05CEF5CEE5CED5CEC5CEB5CEA5CE95CE85CE75CE65CE55CE4",
		x"FFFFFFFFFFFFFFFF5CFF5CFE5CFD5CFC5CFB5CFA5CF95CF85CF75CF65CF55CF4",
		x"5D0F5D0E5D0D5D0C5D0B5D0A5D095D085D075D065D055D045D035D025D015D00",
		x"5D1F5D1E5D1D5D1C5D1B5D1A5D195D185D175D165D155D145D135D125D115D10",
		x"5D2F5D2E5D2D5D2C5D2B5D2A5D295D285D275D265D255D245D235D225D215D20",
		x"5D3F5D3E5D3D5D3C5D3B5D3A5D395D385D375D365D355D345D335D325D315D30",
		x"5D4B5D4A5D495D485D475D465D455D445D435D425D415D40FFFFFFFFFFFFFFFF",
		x"5D5B5D5A5D595D585D575D565D555D545D535D525D515D505D4F5D4E5D4D5D4C",
		x"5D6B5D6A5D695D685D675D665D655D645D635D625D615D605D5F5D5E5D5D5D5C",
		x"5D7B5D7A5D795D785D775D765D755D745D735D725D715D705D6F5D6E5D6D5D6C",
		x"5D875D865D855D845D835D825D815D80FFFFFFFFFFFFFFFF5D7F5D7E5D7D5D7C",
		x"5D975D965D955D945D935D925D915D905D8F5D8E5D8D5D8C5D8B5D8A5D895D88",
		x"5DA75DA65DA55DA45DA35DA25DA15DA05D9F5D9E5D9D5D9C5D9B5D9A5D995D98",
		x"5DB75DB65DB55DB45DB35DB25DB15DB05DAF5DAE5DAD5DAC5DAB5DAA5DA95DA8",
		x"5DC35DC25DC15DC0FFFFFFFFFFFFFFFF5DBF5DBE5DBD5DBC5DBB5DBA5DB95DB8",
		x"5DD35DD25DD15DD05DCF5DCE5DCD5DCC5DCB5DCA5DC95DC85DC75DC65DC55DC4",
		x"5DE35DE25DE15DE05DDF5DDE5DDD5DDC5DDB5DDA5DD95DD85DD75DD65DD55DD4",
		x"5DF35DF25DF15DF05DEF5DEE5DED5DEC5DEB5DEA5DE95DE85DE75DE65DE55DE4",
		x"FFFFFFFFFFFFFFFF5DFF5DFE5DFD5DFC5DFB5DFA5DF95DF85DF75DF65DF55DF4",
		x"5E0F5E0E5E0D5E0C5E0B5E0A5E095E085E075E065E055E045E035E025E015E00",
		x"5E1F5E1E5E1D5E1C5E1B5E1A5E195E185E175E165E155E145E135E125E115E10",
		x"5E2F5E2E5E2D5E2C5E2B5E2A5E295E285E275E265E255E245E235E225E215E20",
		x"5E3F5E3E5E3D5E3C5E3B5E3A5E395E385E375E365E355E345E335E325E315E30",
		x"5E4B5E4A5E495E485E475E465E455E445E435E425E415E40FFFFFFFFFFFFFFFF",
		x"5E5B5E5A5E595E585E575E565E555E545E535E525E515E505E4F5E4E5E4D5E4C",
		x"5E6B5E6A5E695E685E675E665E655E645E635E625E615E605E5F5E5E5E5D5E5C",
		x"5E7B5E7A5E795E785E775E765E755E745E735E725E715E705E6F5E6E5E6D5E6C",
		x"5E875E865E855E845E835E825E815E80FFFFFFFFFFFFFFFF5E7F5E7E5E7D5E7C",
		x"5E975E965E955E945E935E925E915E905E8F5E8E5E8D5E8C5E8B5E8A5E895E88",
		x"5EA75EA65EA55EA45EA35EA25EA15EA05E9F5E9E5E9D5E9C5E9B5E9A5E995E98",
		x"5EB75EB65EB55EB45EB35EB25EB15EB05EAF5EAE5EAD5EAC5EAB5EAA5EA95EA8",
		x"5EC35EC25EC15EC0FFFFFFFFFFFFFFFF5EBF5EBE5EBD5EBC5EBB5EBA5EB95EB8",
		x"5ED35ED25ED15ED05ECF5ECE5ECD5ECC5ECB5ECA5EC95EC85EC75EC65EC55EC4",
		x"5EE35EE25EE15EE05EDF5EDE5EDD5EDC5EDB5EDA5ED95ED85ED75ED65ED55ED4",
		x"5EF35EF25EF15EF05EEF5EEE5EED5EEC5EEB5EEA5EE95EE85EE75EE65EE55EE4",
		x"FFFFFFFFFFFFFFFF5EFF5EFE5EFD5EFC5EFB5EFA5EF95EF85EF75EF65EF55EF4",
		x"5F0F5F0E5F0D5F0C5F0B5F0A5F095F085F075F065F055F045F035F025F015F00",
		x"5F1F5F1E5F1D5F1C5F1B5F1A5F195F185F175F165F155F145F135F125F115F10",
		x"5F2F5F2E5F2D5F2C5F2B5F2A5F295F285F275F265F255F245F235F225F215F20",
		x"5F3F5F3E5F3D5F3C5F3B5F3A5F395F385F375F365F355F345F335F325F315F30",
		x"5F4B5F4A5F495F485F475F465F455F445F435F425F415F40FFFFFFFFFFFFFFFF",
		x"5F5B5F5A5F595F585F575F565F555F545F535F525F515F505F4F5F4E5F4D5F4C",
		x"5F6B5F6A5F695F685F675F665F655F645F635F625F615F605F5F5F5E5F5D5F5C",
		x"5F7B5F7A5F795F785F775F765F755F745F735F725F715F705F6F5F6E5F6D5F6C",
		x"5F875F865F855F845F835F825F815F80FFFFFFFFFFFFFFFF5F7F5F7E5F7D5F7C",
		x"5F975F965F955F945F935F925F915F905F8F5F8E5F8D5F8C5F8B5F8A5F895F88",
		x"5FA75FA65FA55FA45FA35FA25FA15FA05F9F5F9E5F9D5F9C5F9B5F9A5F995F98",
		x"5FB75FB65FB55FB45FB35FB25FB15FB05FAF5FAE5FAD5FAC5FAB5FAA5FA95FA8",
		x"5FC35FC25FC15FC0FFFFFFFFFFFFFFFF5FBF5FBE5FBD5FBC5FBB5FBA5FB95FB8",
		x"5FD35FD25FD15FD05FCF5FCE5FCD5FCC5FCB5FCA5FC95FC85FC75FC65FC55FC4",
		x"5FE35FE25FE15FE05FDF5FDE5FDD5FDC5FDB5FDA5FD95FD85FD75FD65FD55FD4",
		x"5FF35FF25FF15FF05FEF5FEE5FED5FEC5FEB5FEA5FE95FE85FE75FE65FE55FE4",
		x"FFFFFFFFFFFFFFFF5FFF5FFE5FFD5FFC5FFB5FFA5FF95FF85FF75FF65FF55FF4",
		x"600F600E600D600C600B600A6009600860076006600560046003600260016000",
		x"601F601E601D601C601B601A6019601860176016601560146013601260116010",
		x"602F602E602D602C602B602A6029602860276026602560246023602260216020",
		x"603F603E603D603C603B603A6039603860376036603560346033603260316030",
		x"604B604A6049604860476046604560446043604260416040FFFFFFFFFFFFFFFF",
		x"605B605A6059605860576056605560546053605260516050604F604E604D604C",
		x"606B606A6069606860676066606560646063606260616060605F605E605D605C",
		x"607B607A6079607860776076607560746073607260716070606F606E606D606C",
		x"60876086608560846083608260816080FFFFFFFFFFFFFFFF607F607E607D607C",
		x"60976096609560946093609260916090608F608E608D608C608B608A60896088",
		x"60A760A660A560A460A360A260A160A0609F609E609D609C609B609A60996098",
		x"60B760B660B560B460B360B260B160B060AF60AE60AD60AC60AB60AA60A960A8",
		x"60C360C260C160C0FFFFFFFFFFFFFFFF60BF60BE60BD60BC60BB60BA60B960B8",
		x"60D360D260D160D060CF60CE60CD60CC60CB60CA60C960C860C760C660C560C4",
		x"60E360E260E160E060DF60DE60DD60DC60DB60DA60D960D860D760D660D560D4",
		x"60F360F260F160F060EF60EE60ED60EC60EB60EA60E960E860E760E660E560E4",
		x"FFFFFFFFFFFFFFFF60FF60FE60FD60FC60FB60FA60F960F860F760F660F560F4",
		x"610F610E610D610C610B610A6109610861076106610561046103610261016100",
		x"611F611E611D611C611B611A6119611861176116611561146113611261116110",
		x"612F612E612D612C612B612A6129612861276126612561246123612261216120",
		x"613F613E613D613C613B613A6139613861376136613561346133613261316130",
		x"614B614A6149614861476146614561446143614261416140FFFFFFFFFFFFFFFF",
		x"615B615A6159615861576156615561546153615261516150614F614E614D614C",
		x"616B616A6169616861676166616561646163616261616160615F615E615D615C",
		x"617B617A6179617861776176617561746173617261716170616F616E616D616C",
		x"61876186618561846183618261816180FFFFFFFFFFFFFFFF617F617E617D617C",
		x"61976196619561946193619261916190618F618E618D618C618B618A61896188",
		x"61A761A661A561A461A361A261A161A0619F619E619D619C619B619A61996198",
		x"61B761B661B561B461B361B261B161B061AF61AE61AD61AC61AB61AA61A961A8",
		x"61C361C261C161C0FFFFFFFFFFFFFFFF61BF61BE61BD61BC61BB61BA61B961B8",
		x"61D361D261D161D061CF61CE61CD61CC61CB61CA61C961C861C761C661C561C4",
		x"61E361E261E161E061DF61DE61DD61DC61DB61DA61D961D861D761D661D561D4",
		x"61F361F261F161F061EF61EE61ED61EC61EB61EA61E961E861E761E661E561E4",
		x"FFFFFFFFFFFFFFFF61FF61FE61FD61FC61FB61FA61F961F861F761F661F561F4",
		x"620F620E620D620C620B620A6209620862076206620562046203620262016200",
		x"621F621E621D621C621B621A6219621862176216621562146213621262116210",
		x"622F622E622D622C622B622A6229622862276226622562246223622262216220",
		x"623F623E623D623C623B623A6239623862376236623562346233623262316230",
		x"624B624A6249624862476246624562446243624262416240FFFFFFFFFFFFFFFF",
		x"625B625A6259625862576256625562546253625262516250624F624E624D624C",
		x"626B626A6269626862676266626562646263626262616260625F625E625D625C",
		x"627B627A6279627862776276627562746273627262716270626F626E626D626C",
		x"62876286628562846283628262816280FFFFFFFFFFFFFFFF627F627E627D627C",
		x"62976296629562946293629262916290628F628E628D628C628B628A62896288",
		x"62A762A662A562A462A362A262A162A0629F629E629D629C629B629A62996298",
		x"62B762B662B562B462B362B262B162B062AF62AE62AD62AC62AB62AA62A962A8",
		x"62C362C262C162C0FFFFFFFFFFFFFFFF62BF62BE62BD62BC62BB62BA62B962B8",
		x"62D362D262D162D062CF62CE62CD62CC62CB62CA62C962C862C762C662C562C4",
		x"62E362E262E162E062DF62DE62DD62DC62DB62DA62D962D862D762D662D562D4",
		x"62F362F262F162F062EF62EE62ED62EC62EB62EA62E962E862E762E662E562E4",
		x"FFFFFFFFFFFFFFFF62FF62FE62FD62FC62FB62FA62F962F862F762F662F562F4",
		x"630F630E630D630C630B630A6309630863076306630563046303630263016300",
		x"631F631E631D631C631B631A6319631863176316631563146313631263116310",
		x"632F632E632D632C632B632A6329632863276326632563246323632263216320",
		x"633F633E633D633C633B633A6339633863376336633563346333633263316330",
		x"634B634A6349634863476346634563446343634263416340FFFFFFFFFFFFFFFF",
		x"635B635A6359635863576356635563546353635263516350634F634E634D634C",
		x"636B636A6369636863676366636563646363636263616360635F635E635D635C",
		x"637B637A6379637863776376637563746373637263716370636F636E636D636C",
		x"63876386638563846383638263816380FFFFFFFFFFFFFFFF637F637E637D637C",
		x"63976396639563946393639263916390638F638E638D638C638B638A63896388",
		x"63A763A663A563A463A363A263A163A0639F639E639D639C639B639A63996398",
		x"63B763B663B563B463B363B263B163B063AF63AE63AD63AC63AB63AA63A963A8",
		x"63C363C263C163C0FFFFFFFFFFFFFFFF63BF63BE63BD63BC63BB63BA63B963B8",
		x"63D363D263D163D063CF63CE63CD63CC63CB63CA63C963C863C763C663C563C4",
		x"63E363E263E163E063DF63DE63DD63DC63DB63DA63D963D863D763D663D563D4",
		x"63F363F263F163F063EF63EE63ED63EC63EB63EA63E963E863E763E663E563E4",
		x"FFFFFFFFFFFFFFFF63FF63FE63FD63FC63FB63FA63F963F863F763F663F563F4",
		x"640F640E640D640C640B640A6409640864076406640564046403640264016400",
		x"641F641E641D641C641B641A6419641864176416641564146413641264116410",
		x"642F642E642D642C642B642A6429642864276426642564246423642264216420",
		x"643F643E643D643C643B643A6439643864376436643564346433643264316430",
		x"644B644A6449644864476446644564446443644264416440FFFFFFFFFFFFFFFF",
		x"645B645A6459645864576456645564546453645264516450644F644E644D644C",
		x"646B646A6469646864676466646564646463646264616460645F645E645D645C",
		x"647B647A6479647864776476647564746473647264716470646F646E646D646C",
		x"64876486648564846483648264816480FFFFFFFFFFFFFFFF647F647E647D647C",
		x"64976496649564946493649264916490648F648E648D648C648B648A64896488",
		x"64A764A664A564A464A364A264A164A0649F649E649D649C649B649A64996498",
		x"64B764B664B564B464B364B264B164B064AF64AE64AD64AC64AB64AA64A964A8",
		x"64C364C264C164C0FFFFFFFFFFFFFFFF64BF64BE64BD64BC64BB64BA64B964B8",
		x"64D364D264D164D064CF64CE64CD64CC64CB64CA64C964C864C764C664C564C4",
		x"64E364E264E164E064DF64DE64DD64DC64DB64DA64D964D864D764D664D564D4",
		x"64F364F264F164F064EF64EE64ED64EC64EB64EA64E964E864E764E664E564E4",
		x"FFFFFFFFFFFFFFFF64FF64FE64FD64FC64FB64FA64F964F864F764F664F564F4",
		x"650F650E650D650C650B650A6509650865076506650565046503650265016500",
		x"651F651E651D651C651B651A6519651865176516651565146513651265116510",
		x"652F652E652D652C652B652A6529652865276526652565246523652265216520",
		x"653F653E653D653C653B653A6539653865376536653565346533653265316530",
		x"654B654A6549654865476546654565446543654265416540FFFFFFFFFFFFFFFF",
		x"655B655A6559655865576556655565546553655265516550654F654E654D654C",
		x"656B656A6569656865676566656565646563656265616560655F655E655D655C",
		x"657B657A6579657865776576657565746573657265716570656F656E656D656C",
		x"65876586658565846583658265816580FFFFFFFFFFFFFFFF657F657E657D657C",
		x"65976596659565946593659265916590658F658E658D658C658B658A65896588",
		x"65A765A665A565A465A365A265A165A0659F659E659D659C659B659A65996598",
		x"65B765B665B565B465B365B265B165B065AF65AE65AD65AC65AB65AA65A965A8",
		x"65C365C265C165C0FFFFFFFFFFFFFFFF65BF65BE65BD65BC65BB65BA65B965B8",
		x"65D365D265D165D065CF65CE65CD65CC65CB65CA65C965C865C765C665C565C4",
		x"65E365E265E165E065DF65DE65DD65DC65DB65DA65D965D865D765D665D565D4",
		x"65F365F265F165F065EF65EE65ED65EC65EB65EA65E965E865E765E665E565E4",
		x"FFFFFFFFFFFFFFFF65FF65FE65FD65FC65FB65FA65F965F865F765F665F565F4",
		x"660F660E660D660C660B660A6609660866076606660566046603660266016600",
		x"661F661E661D661C661B661A6619661866176616661566146613661266116610",
		x"662F662E662D662C662B662A6629662866276626662566246623662266216620",
		x"663F663E663D663C663B663A6639663866376636663566346633663266316630",
		x"664B664A6649664866476646664566446643664266416640FFFFFFFFFFFFFFFF",
		x"665B665A6659665866576656665566546653665266516650664F664E664D664C",
		x"666B666A6669666866676666666566646663666266616660665F665E665D665C",
		x"667B667A6679667866776676667566746673667266716670666F666E666D666C",
		x"66876686668566846683668266816680FFFFFFFFFFFFFFFF667F667E667D667C",
		x"66976696669566946693669266916690668F668E668D668C668B668A66896688",
		x"66A766A666A566A466A366A266A166A0669F669E669D669C669B669A66996698",
		x"66B766B666B566B466B366B266B166B066AF66AE66AD66AC66AB66AA66A966A8",
		x"66C366C266C166C0FFFFFFFFFFFFFFFF66BF66BE66BD66BC66BB66BA66B966B8",
		x"66D366D266D166D066CF66CE66CD66CC66CB66CA66C966C866C766C666C566C4",
		x"66E366E266E166E066DF66DE66DD66DC66DB66DA66D966D866D766D666D566D4",
		x"66F366F266F166F066EF66EE66ED66EC66EB66EA66E966E866E766E666E566E4",
		x"FFFFFFFFFFFFFFFF66FF66FE66FD66FC66FB66FA66F966F866F766F666F566F4",
		x"670F670E670D670C670B670A6709670867076706670567046703670267016700",
		x"671F671E671D671C671B671A6719671867176716671567146713671267116710",
		x"672F672E672D672C672B672A6729672867276726672567246723672267216720",
		x"673F673E673D673C673B673A6739673867376736673567346733673267316730",
		x"674B674A6749674867476746674567446743674267416740FFFFFFFFFFFFFFFF",
		x"675B675A6759675867576756675567546753675267516750674F674E674D674C",
		x"676B676A6769676867676766676567646763676267616760675F675E675D675C",
		x"677B677A6779677867776776677567746773677267716770676F676E676D676C",
		x"67876786678567846783678267816780FFFFFFFFFFFFFFFF677F677E677D677C",
		x"67976796679567946793679267916790678F678E678D678C678B678A67896788",
		x"67A767A667A567A467A367A267A167A0679F679E679D679C679B679A67996798",
		x"67B767B667B567B467B367B267B167B067AF67AE67AD67AC67AB67AA67A967A8",
		x"67C367C267C167C0FFFFFFFFFFFFFFFF67BF67BE67BD67BC67BB67BA67B967B8",
		x"67D367D267D167D067CF67CE67CD67CC67CB67CA67C967C867C767C667C567C4",
		x"67E367E267E167E067DF67DE67DD67DC67DB67DA67D967D867D767D667D567D4",
		x"67F367F267F167F067EF67EE67ED67EC67EB67EA67E967E867E767E667E567E4",
		x"FFFFFFFFFFFFFFFF67FF67FE67FD67FC67FB67FA67F967F867F767F667F567F4",
		x"680F680E680D680C680B680A6809680868076806680568046803680268016800",
		x"681F681E681D681C681B681A6819681868176816681568146813681268116810",
		x"682F682E682D682C682B682A6829682868276826682568246823682268216820",
		x"683F683E683D683C683B683A6839683868376836683568346833683268316830",
		x"684B684A6849684868476846684568446843684268416840FFFFFFFFFFFFFFFF",
		x"685B685A6859685868576856685568546853685268516850684F684E684D684C",
		x"686B686A6869686868676866686568646863686268616860685F685E685D685C",
		x"687B687A6879687868776876687568746873687268716870686F686E686D686C",
		x"68876886688568846883688268816880FFFFFFFFFFFFFFFF687F687E687D687C",
		x"68976896689568946893689268916890688F688E688D688C688B688A68896888",
		x"68A768A668A568A468A368A268A168A0689F689E689D689C689B689A68996898",
		x"68B768B668B568B468B368B268B168B068AF68AE68AD68AC68AB68AA68A968A8",
		x"68C368C268C168C0FFFFFFFFFFFFFFFF68BF68BE68BD68BC68BB68BA68B968B8",
		x"68D368D268D168D068CF68CE68CD68CC68CB68CA68C968C868C768C668C568C4",
		x"68E368E268E168E068DF68DE68DD68DC68DB68DA68D968D868D768D668D568D4",
		x"68F368F268F168F068EF68EE68ED68EC68EB68EA68E968E868E768E668E568E4",
		x"FFFFFFFFFFFFFFFF68FF68FE68FD68FC68FB68FA68F968F868F768F668F568F4",
		x"690F690E690D690C690B690A6909690869076906690569046903690269016900",
		x"691F691E691D691C691B691A6919691869176916691569146913691269116910",
		x"692F692E692D692C692B692A6929692869276926692569246923692269216920",
		x"693F693E693D693C693B693A6939693869376936693569346933693269316930",
		x"694B694A6949694869476946694569446943694269416940FFFFFFFFFFFFFFFF",
		x"695B695A6959695869576956695569546953695269516950694F694E694D694C",
		x"696B696A6969696869676966696569646963696269616960695F695E695D695C",
		x"697B697A6979697869776976697569746973697269716970696F696E696D696C",
		x"69876986698569846983698269816980FFFFFFFFFFFFFFFF697F697E697D697C",
		x"69976996699569946993699269916990698F698E698D698C698B698A69896988",
		x"69A769A669A569A469A369A269A169A0699F699E699D699C699B699A69996998",
		x"69B769B669B569B469B369B269B169B069AF69AE69AD69AC69AB69AA69A969A8",
		x"69C369C269C169C0FFFFFFFFFFFFFFFF69BF69BE69BD69BC69BB69BA69B969B8",
		x"69D369D269D169D069CF69CE69CD69CC69CB69CA69C969C869C769C669C569C4",
		x"69E369E269E169E069DF69DE69DD69DC69DB69DA69D969D869D769D669D569D4",
		x"69F369F269F169F069EF69EE69ED69EC69EB69EA69E969E869E769E669E569E4",
		x"FFFFFFFFFFFFFFFF69FF69FE69FD69FC69FB69FA69F969F869F769F669F569F4",
		x"6A0F6A0E6A0D6A0C6A0B6A0A6A096A086A076A066A056A046A036A026A016A00",
		x"6A1F6A1E6A1D6A1C6A1B6A1A6A196A186A176A166A156A146A136A126A116A10",
		x"6A2F6A2E6A2D6A2C6A2B6A2A6A296A286A276A266A256A246A236A226A216A20",
		x"6A3F6A3E6A3D6A3C6A3B6A3A6A396A386A376A366A356A346A336A326A316A30",
		x"6A4B6A4A6A496A486A476A466A456A446A436A426A416A40FFFFFFFFFFFFFFFF",
		x"6A5B6A5A6A596A586A576A566A556A546A536A526A516A506A4F6A4E6A4D6A4C",
		x"6A6B6A6A6A696A686A676A666A656A646A636A626A616A606A5F6A5E6A5D6A5C",
		x"6A7B6A7A6A796A786A776A766A756A746A736A726A716A706A6F6A6E6A6D6A6C",
		x"6A876A866A856A846A836A826A816A80FFFFFFFFFFFFFFFF6A7F6A7E6A7D6A7C",
		x"6A976A966A956A946A936A926A916A906A8F6A8E6A8D6A8C6A8B6A8A6A896A88",
		x"6AA76AA66AA56AA46AA36AA26AA16AA06A9F6A9E6A9D6A9C6A9B6A9A6A996A98",
		x"6AB76AB66AB56AB46AB36AB26AB16AB06AAF6AAE6AAD6AAC6AAB6AAA6AA96AA8",
		x"6AC36AC26AC16AC0FFFFFFFFFFFFFFFF6ABF6ABE6ABD6ABC6ABB6ABA6AB96AB8",
		x"6AD36AD26AD16AD06ACF6ACE6ACD6ACC6ACB6ACA6AC96AC86AC76AC66AC56AC4",
		x"6AE36AE26AE16AE06ADF6ADE6ADD6ADC6ADB6ADA6AD96AD86AD76AD66AD56AD4",
		x"6AF36AF26AF16AF06AEF6AEE6AED6AEC6AEB6AEA6AE96AE86AE76AE66AE56AE4",
		x"FFFFFFFFFFFFFFFF6AFF6AFE6AFD6AFC6AFB6AFA6AF96AF86AF76AF66AF56AF4",
		x"6B0F6B0E6B0D6B0C6B0B6B0A6B096B086B076B066B056B046B036B026B016B00",
		x"6B1F6B1E6B1D6B1C6B1B6B1A6B196B186B176B166B156B146B136B126B116B10",
		x"6B2F6B2E6B2D6B2C6B2B6B2A6B296B286B276B266B256B246B236B226B216B20",
		x"6B3F6B3E6B3D6B3C6B3B6B3A6B396B386B376B366B356B346B336B326B316B30",
		x"6B4B6B4A6B496B486B476B466B456B446B436B426B416B40FFFFFFFFFFFFFFFF",
		x"6B5B6B5A6B596B586B576B566B556B546B536B526B516B506B4F6B4E6B4D6B4C",
		x"6B6B6B6A6B696B686B676B666B656B646B636B626B616B606B5F6B5E6B5D6B5C",
		x"6B7B6B7A6B796B786B776B766B756B746B736B726B716B706B6F6B6E6B6D6B6C",
		x"6B876B866B856B846B836B826B816B80FFFFFFFFFFFFFFFF6B7F6B7E6B7D6B7C",
		x"6B976B966B956B946B936B926B916B906B8F6B8E6B8D6B8C6B8B6B8A6B896B88",
		x"6BA76BA66BA56BA46BA36BA26BA16BA06B9F6B9E6B9D6B9C6B9B6B9A6B996B98",
		x"6BB76BB66BB56BB46BB36BB26BB16BB06BAF6BAE6BAD6BAC6BAB6BAA6BA96BA8",
		x"6BC36BC26BC16BC0FFFFFFFFFFFFFFFF6BBF6BBE6BBD6BBC6BBB6BBA6BB96BB8",
		x"6BD36BD26BD16BD06BCF6BCE6BCD6BCC6BCB6BCA6BC96BC86BC76BC66BC56BC4",
		x"6BE36BE26BE16BE06BDF6BDE6BDD6BDC6BDB6BDA6BD96BD86BD76BD66BD56BD4",
		x"6BF36BF26BF16BF06BEF6BEE6BED6BEC6BEB6BEA6BE96BE86BE76BE66BE56BE4",
		x"FFFFFFFFFFFFFFFF6BFF6BFE6BFD6BFC6BFB6BFA6BF96BF86BF76BF66BF56BF4",
		x"6C0F6C0E6C0D6C0C6C0B6C0A6C096C086C076C066C056C046C036C026C016C00",
		x"6C1F6C1E6C1D6C1C6C1B6C1A6C196C186C176C166C156C146C136C126C116C10",
		x"6C2F6C2E6C2D6C2C6C2B6C2A6C296C286C276C266C256C246C236C226C216C20",
		x"6C3F6C3E6C3D6C3C6C3B6C3A6C396C386C376C366C356C346C336C326C316C30",
		x"6C4B6C4A6C496C486C476C466C456C446C436C426C416C40FFFFFFFFFFFFFFFF",
		x"6C5B6C5A6C596C586C576C566C556C546C536C526C516C506C4F6C4E6C4D6C4C",
		x"6C6B6C6A6C696C686C676C666C656C646C636C626C616C606C5F6C5E6C5D6C5C",
		x"6C7B6C7A6C796C786C776C766C756C746C736C726C716C706C6F6C6E6C6D6C6C",
		x"6C876C866C856C846C836C826C816C80FFFFFFFFFFFFFFFF6C7F6C7E6C7D6C7C",
		x"6C976C966C956C946C936C926C916C906C8F6C8E6C8D6C8C6C8B6C8A6C896C88",
		x"6CA76CA66CA56CA46CA36CA26CA16CA06C9F6C9E6C9D6C9C6C9B6C9A6C996C98",
		x"6CB76CB66CB56CB46CB36CB26CB16CB06CAF6CAE6CAD6CAC6CAB6CAA6CA96CA8",
		x"6CC36CC26CC16CC0FFFFFFFFFFFFFFFF6CBF6CBE6CBD6CBC6CBB6CBA6CB96CB8",
		x"6CD36CD26CD16CD06CCF6CCE6CCD6CCC6CCB6CCA6CC96CC86CC76CC66CC56CC4",
		x"6CE36CE26CE16CE06CDF6CDE6CDD6CDC6CDB6CDA6CD96CD86CD76CD66CD56CD4",
		x"6CF36CF26CF16CF06CEF6CEE6CED6CEC6CEB6CEA6CE96CE86CE76CE66CE56CE4",
		x"FFFFFFFFFFFFFFFF6CFF6CFE6CFD6CFC6CFB6CFA6CF96CF86CF76CF66CF56CF4",
		x"6D0F6D0E6D0D6D0C6D0B6D0A6D096D086D076D066D056D046D036D026D016D00",
		x"6D1F6D1E6D1D6D1C6D1B6D1A6D196D186D176D166D156D146D136D126D116D10",
		x"6D2F6D2E6D2D6D2C6D2B6D2A6D296D286D276D266D256D246D236D226D216D20",
		x"6D3F6D3E6D3D6D3C6D3B6D3A6D396D386D376D366D356D346D336D326D316D30",
		x"6D4B6D4A6D496D486D476D466D456D446D436D426D416D40FFFFFFFFFFFFFFFF",
		x"6D5B6D5A6D596D586D576D566D556D546D536D526D516D506D4F6D4E6D4D6D4C",
		x"6D6B6D6A6D696D686D676D666D656D646D636D626D616D606D5F6D5E6D5D6D5C",
		x"6D7B6D7A6D796D786D776D766D756D746D736D726D716D706D6F6D6E6D6D6D6C",
		x"6D876D866D856D846D836D826D816D80FFFFFFFFFFFFFFFF6D7F6D7E6D7D6D7C",
		x"6D976D966D956D946D936D926D916D906D8F6D8E6D8D6D8C6D8B6D8A6D896D88",
		x"6DA76DA66DA56DA46DA36DA26DA16DA06D9F6D9E6D9D6D9C6D9B6D9A6D996D98",
		x"6DB76DB66DB56DB46DB36DB26DB16DB06DAF6DAE6DAD6DAC6DAB6DAA6DA96DA8",
		x"6DC36DC26DC16DC0FFFFFFFFFFFFFFFF6DBF6DBE6DBD6DBC6DBB6DBA6DB96DB8",
		x"6DD36DD26DD16DD06DCF6DCE6DCD6DCC6DCB6DCA6DC96DC86DC76DC66DC56DC4",
		x"6DE36DE26DE16DE06DDF6DDE6DDD6DDC6DDB6DDA6DD96DD86DD76DD66DD56DD4",
		x"6DF36DF26DF16DF06DEF6DEE6DED6DEC6DEB6DEA6DE96DE86DE76DE66DE56DE4",
		x"FFFFFFFFFFFFFFFF6DFF6DFE6DFD6DFC6DFB6DFA6DF96DF86DF76DF66DF56DF4",
		x"6E0F6E0E6E0D6E0C6E0B6E0A6E096E086E076E066E056E046E036E026E016E00",
		x"6E1F6E1E6E1D6E1C6E1B6E1A6E196E186E176E166E156E146E136E126E116E10",
		x"6E2F6E2E6E2D6E2C6E2B6E2A6E296E286E276E266E256E246E236E226E216E20",
		x"6E3F6E3E6E3D6E3C6E3B6E3A6E396E386E376E366E356E346E336E326E316E30",
		x"6E4B6E4A6E496E486E476E466E456E446E436E426E416E40FFFFFFFFFFFFFFFF",
		x"6E5B6E5A6E596E586E576E566E556E546E536E526E516E506E4F6E4E6E4D6E4C",
		x"6E6B6E6A6E696E686E676E666E656E646E636E626E616E606E5F6E5E6E5D6E5C",
		x"6E7B6E7A6E796E786E776E766E756E746E736E726E716E706E6F6E6E6E6D6E6C",
		x"6E876E866E856E846E836E826E816E80FFFFFFFFFFFFFFFF6E7F6E7E6E7D6E7C",
		x"6E976E966E956E946E936E926E916E906E8F6E8E6E8D6E8C6E8B6E8A6E896E88",
		x"6EA76EA66EA56EA46EA36EA26EA16EA06E9F6E9E6E9D6E9C6E9B6E9A6E996E98",
		x"6EB76EB66EB56EB46EB36EB26EB16EB06EAF6EAE6EAD6EAC6EAB6EAA6EA96EA8",
		x"6EC36EC26EC16EC0FFFFFFFFFFFFFFFF6EBF6EBE6EBD6EBC6EBB6EBA6EB96EB8",
		x"6ED36ED26ED16ED06ECF6ECE6ECD6ECC6ECB6ECA6EC96EC86EC76EC66EC56EC4",
		x"6EE36EE26EE16EE06EDF6EDE6EDD6EDC6EDB6EDA6ED96ED86ED76ED66ED56ED4",
		x"6EF36EF26EF16EF06EEF6EEE6EED6EEC6EEB6EEA6EE96EE86EE76EE66EE56EE4",
		x"FFFFFFFFFFFFFFFF6EFF6EFE6EFD6EFC6EFB6EFA6EF96EF86EF76EF66EF56EF4",
		x"6F0F6F0E6F0D6F0C6F0B6F0A6F096F086F076F066F056F046F036F026F016F00",
		x"6F1F6F1E6F1D6F1C6F1B6F1A6F196F186F176F166F156F146F136F126F116F10",
		x"6F2F6F2E6F2D6F2C6F2B6F2A6F296F286F276F266F256F246F236F226F216F20",
		x"6F3F6F3E6F3D6F3C6F3B6F3A6F396F386F376F366F356F346F336F326F316F30",
		x"6F4B6F4A6F496F486F476F466F456F446F436F426F416F40FFFFFFFFFFFFFFFF",
		x"6F5B6F5A6F596F586F576F566F556F546F536F526F516F506F4F6F4E6F4D6F4C",
		x"6F6B6F6A6F696F686F676F666F656F646F636F626F616F606F5F6F5E6F5D6F5C",
		x"6F7B6F7A6F796F786F776F766F756F746F736F726F716F706F6F6F6E6F6D6F6C",
		x"6F876F866F856F846F836F826F816F80FFFFFFFFFFFFFFFF6F7F6F7E6F7D6F7C",
		x"6F976F966F956F946F936F926F916F906F8F6F8E6F8D6F8C6F8B6F8A6F896F88",
		x"6FA76FA66FA56FA46FA36FA26FA16FA06F9F6F9E6F9D6F9C6F9B6F9A6F996F98",
		x"6FB76FB66FB56FB46FB36FB26FB16FB06FAF6FAE6FAD6FAC6FAB6FAA6FA96FA8",
		x"6FC36FC26FC16FC0FFFFFFFFFFFFFFFF6FBF6FBE6FBD6FBC6FBB6FBA6FB96FB8",
		x"6FD36FD26FD16FD06FCF6FCE6FCD6FCC6FCB6FCA6FC96FC86FC76FC66FC56FC4",
		x"6FE36FE26FE16FE06FDF6FDE6FDD6FDC6FDB6FDA6FD96FD86FD76FD66FD56FD4",
		x"6FF36FF26FF16FF06FEF6FEE6FED6FEC6FEB6FEA6FE96FE86FE76FE66FE56FE4",
		x"FFFFFFFFFFFFFFFF6FFF6FFE6FFD6FFC6FFB6FFA6FF96FF86FF76FF66FF56FF4",
		x"700F700E700D700C700B700A7009700870077006700570047003700270017000",
		x"701F701E701D701C701B701A7019701870177016701570147013701270117010",
		x"702F702E702D702C702B702A7029702870277026702570247023702270217020",
		x"703F703E703D703C703B703A7039703870377036703570347033703270317030",
		x"704B704A7049704870477046704570447043704270417040FFFFFFFFFFFFFFFF",
		x"705B705A7059705870577056705570547053705270517050704F704E704D704C",
		x"706B706A7069706870677066706570647063706270617060705F705E705D705C",
		x"707B707A7079707870777076707570747073707270717070706F706E706D706C",
		x"70877086708570847083708270817080FFFFFFFFFFFFFFFF707F707E707D707C",
		x"70977096709570947093709270917090708F708E708D708C708B708A70897088",
		x"70A770A670A570A470A370A270A170A0709F709E709D709C709B709A70997098",
		x"70B770B670B570B470B370B270B170B070AF70AE70AD70AC70AB70AA70A970A8",
		x"70C370C270C170C0FFFFFFFFFFFFFFFF70BF70BE70BD70BC70BB70BA70B970B8",
		x"70D370D270D170D070CF70CE70CD70CC70CB70CA70C970C870C770C670C570C4",
		x"70E370E270E170E070DF70DE70DD70DC70DB70DA70D970D870D770D670D570D4",
		x"70F370F270F170F070EF70EE70ED70EC70EB70EA70E970E870E770E670E570E4",
		x"FFFFFFFFFFFFFFFF70FF70FE70FD70FC70FB70FA70F970F870F770F670F570F4",
		x"710F710E710D710C710B710A7109710871077106710571047103710271017100",
		x"711F711E711D711C711B711A7119711871177116711571147113711271117110",
		x"712F712E712D712C712B712A7129712871277126712571247123712271217120",
		x"713F713E713D713C713B713A7139713871377136713571347133713271317130",
		x"714B714A7149714871477146714571447143714271417140FFFFFFFFFFFFFFFF",
		x"715B715A7159715871577156715571547153715271517150714F714E714D714C",
		x"716B716A7169716871677166716571647163716271617160715F715E715D715C",
		x"717B717A7179717871777176717571747173717271717170716F716E716D716C",
		x"71877186718571847183718271817180FFFFFFFFFFFFFFFF717F717E717D717C",
		x"71977196719571947193719271917190718F718E718D718C718B718A71897188",
		x"71A771A671A571A471A371A271A171A0719F719E719D719C719B719A71997198",
		x"71B771B671B571B471B371B271B171B071AF71AE71AD71AC71AB71AA71A971A8",
		x"71C371C271C171C0FFFFFFFFFFFFFFFF71BF71BE71BD71BC71BB71BA71B971B8",
		x"71D371D271D171D071CF71CE71CD71CC71CB71CA71C971C871C771C671C571C4",
		x"71E371E271E171E071DF71DE71DD71DC71DB71DA71D971D871D771D671D571D4",
		x"71F371F271F171F071EF71EE71ED71EC71EB71EA71E971E871E771E671E571E4",
		x"FFFFFFFFFFFFFFFF71FF71FE71FD71FC71FB71FA71F971F871F771F671F571F4",
		x"720F720E720D720C720B720A7209720872077206720572047203720272017200",
		x"721F721E721D721C721B721A7219721872177216721572147213721272117210",
		x"722F722E722D722C722B722A7229722872277226722572247223722272217220",
		x"723F723E723D723C723B723A7239723872377236723572347233723272317230",
		x"724B724A7249724872477246724572447243724272417240FFFFFFFFFFFFFFFF",
		x"725B725A7259725872577256725572547253725272517250724F724E724D724C",
		x"726B726A7269726872677266726572647263726272617260725F725E725D725C",
		x"727B727A7279727872777276727572747273727272717270726F726E726D726C",
		x"72877286728572847283728272817280FFFFFFFFFFFFFFFF727F727E727D727C",
		x"72977296729572947293729272917290728F728E728D728C728B728A72897288",
		x"72A772A672A572A472A372A272A172A0729F729E729D729C729B729A72997298",
		x"72B772B672B572B472B372B272B172B072AF72AE72AD72AC72AB72AA72A972A8",
		x"72C372C272C172C0FFFFFFFFFFFFFFFF72BF72BE72BD72BC72BB72BA72B972B8",
		x"72D372D272D172D072CF72CE72CD72CC72CB72CA72C972C872C772C672C572C4",
		x"72E372E272E172E072DF72DE72DD72DC72DB72DA72D972D872D772D672D572D4",
		x"72F372F272F172F072EF72EE72ED72EC72EB72EA72E972E872E772E672E572E4",
		x"FFFFFFFFFFFFFFFF72FF72FE72FD72FC72FB72FA72F972F872F772F672F572F4",
		x"730F730E730D730C730B730A7309730873077306730573047303730273017300",
		x"731F731E731D731C731B731A7319731873177316731573147313731273117310",
		x"732F732E732D732C732B732A7329732873277326732573247323732273217320",
		x"733F733E733D733C733B733A7339733873377336733573347333733273317330",
		x"734B734A7349734873477346734573447343734273417340FFFFFFFFFFFFFFFF",
		x"735B735A7359735873577356735573547353735273517350734F734E734D734C",
		x"736B736A7369736873677366736573647363736273617360735F735E735D735C",
		x"737B737A7379737873777376737573747373737273717370736F736E736D736C",
		x"73877386738573847383738273817380FFFFFFFFFFFFFFFF737F737E737D737C",
		x"73977396739573947393739273917390738F738E738D738C738B738A73897388",
		x"73A773A673A573A473A373A273A173A0739F739E739D739C739B739A73997398",
		x"73B773B673B573B473B373B273B173B073AF73AE73AD73AC73AB73AA73A973A8",
		x"73C373C273C173C0FFFFFFFFFFFFFFFF73BF73BE73BD73BC73BB73BA73B973B8",
		x"73D373D273D173D073CF73CE73CD73CC73CB73CA73C973C873C773C673C573C4",
		x"73E373E273E173E073DF73DE73DD73DC73DB73DA73D973D873D773D673D573D4",
		x"73F373F273F173F073EF73EE73ED73EC73EB73EA73E973E873E773E673E573E4",
		x"FFFFFFFFFFFFFFFF73FF73FE73FD73FC73FB73FA73F973F873F773F673F573F4",
		x"740F740E740D740C740B740A7409740874077406740574047403740274017400",
		x"741F741E741D741C741B741A7419741874177416741574147413741274117410",
		x"742F742E742D742C742B742A7429742874277426742574247423742274217420",
		x"743F743E743D743C743B743A7439743874377436743574347433743274317430",
		x"744B744A7449744874477446744574447443744274417440FFFFFFFFFFFFFFFF",
		x"745B745A7459745874577456745574547453745274517450744F744E744D744C",
		x"746B746A7469746874677466746574647463746274617460745F745E745D745C",
		x"747B747A7479747874777476747574747473747274717470746F746E746D746C",
		x"74877486748574847483748274817480FFFFFFFFFFFFFFFF747F747E747D747C",
		x"74977496749574947493749274917490748F748E748D748C748B748A74897488",
		x"74A774A674A574A474A374A274A174A0749F749E749D749C749B749A74997498",
		x"74B774B674B574B474B374B274B174B074AF74AE74AD74AC74AB74AA74A974A8",
		x"74C374C274C174C0FFFFFFFFFFFFFFFF74BF74BE74BD74BC74BB74BA74B974B8",
		x"74D374D274D174D074CF74CE74CD74CC74CB74CA74C974C874C774C674C574C4",
		x"74E374E274E174E074DF74DE74DD74DC74DB74DA74D974D874D774D674D574D4",
		x"74F374F274F174F074EF74EE74ED74EC74EB74EA74E974E874E774E674E574E4",
		x"FFFFFFFFFFFFFFFF74FF74FE74FD74FC74FB74FA74F974F874F774F674F574F4",
		x"750F750E750D750C750B750A7509750875077506750575047503750275017500",
		x"751F751E751D751C751B751A7519751875177516751575147513751275117510",
		x"752F752E752D752C752B752A7529752875277526752575247523752275217520",
		x"753F753E753D753C753B753A7539753875377536753575347533753275317530",
		x"754B754A7549754875477546754575447543754275417540FFFFFFFFFFFFFFFF",
		x"755B755A7559755875577556755575547553755275517550754F754E754D754C",
		x"756B756A7569756875677566756575647563756275617560755F755E755D755C",
		x"757B757A7579757875777576757575747573757275717570756F756E756D756C",
		x"75877586758575847583758275817580FFFFFFFFFFFFFFFF757F757E757D757C",
		x"75977596759575947593759275917590758F758E758D758C758B758A75897588",
		x"75A775A675A575A475A375A275A175A0759F759E759D759C759B759A75997598",
		x"75B775B675B575B475B375B275B175B075AF75AE75AD75AC75AB75AA75A975A8",
		x"75C375C275C175C0FFFFFFFFFFFFFFFF75BF75BE75BD75BC75BB75BA75B975B8",
		x"75D375D275D175D075CF75CE75CD75CC75CB75CA75C975C875C775C675C575C4",
		x"75E375E275E175E075DF75DE75DD75DC75DB75DA75D975D875D775D675D575D4",
		x"75F375F275F175F075EF75EE75ED75EC75EB75EA75E975E875E775E675E575E4",
		x"FFFFFFFFFFFFFFFF75FF75FE75FD75FC75FB75FA75F975F875F775F675F575F4",
		x"760F760E760D760C760B760A7609760876077606760576047603760276017600",
		x"761F761E761D761C761B761A7619761876177616761576147613761276117610",
		x"762F762E762D762C762B762A7629762876277626762576247623762276217620",
		x"763F763E763D763C763B763A7639763876377636763576347633763276317630",
		x"764B764A7649764876477646764576447643764276417640FFFFFFFFFFFFFFFF",
		x"765B765A7659765876577656765576547653765276517650764F764E764D764C",
		x"766B766A7669766876677666766576647663766276617660765F765E765D765C",
		x"767B767A7679767876777676767576747673767276717670766F766E766D766C",
		x"76877686768576847683768276817680FFFFFFFFFFFFFFFF767F767E767D767C",
		x"76977696769576947693769276917690768F768E768D768C768B768A76897688",
		x"76A776A676A576A476A376A276A176A0769F769E769D769C769B769A76997698",
		x"76B776B676B576B476B376B276B176B076AF76AE76AD76AC76AB76AA76A976A8",
		x"76C376C276C176C0FFFFFFFFFFFFFFFF76BF76BE76BD76BC76BB76BA76B976B8",
		x"76D376D276D176D076CF76CE76CD76CC76CB76CA76C976C876C776C676C576C4",
		x"76E376E276E176E076DF76DE76DD76DC76DB76DA76D976D876D776D676D576D4",
		x"76F376F276F176F076EF76EE76ED76EC76EB76EA76E976E876E776E676E576E4",
		x"FFFFFFFFFFFFFFFF76FF76FE76FD76FC76FB76FA76F976F876F776F676F576F4",
		x"770F770E770D770C770B770A7709770877077706770577047703770277017700",
		x"771F771E771D771C771B771A7719771877177716771577147713771277117710",
		x"772F772E772D772C772B772A7729772877277726772577247723772277217720",
		x"773F773E773D773C773B773A7739773877377736773577347733773277317730",
		x"774B774A7749774877477746774577447743774277417740FFFFFFFFFFFFFFFF",
		x"775B775A7759775877577756775577547753775277517750774F774E774D774C",
		x"776B776A7769776877677766776577647763776277617760775F775E775D775C",
		x"777B777A7779777877777776777577747773777277717770776F776E776D776C",
		x"77877786778577847783778277817780FFFFFFFFFFFFFFFF777F777E777D777C",
		x"77977796779577947793779277917790778F778E778D778C778B778A77897788",
		x"77A777A677A577A477A377A277A177A0779F779E779D779C779B779A77997798",
		x"77B777B677B577B477B377B277B177B077AF77AE77AD77AC77AB77AA77A977A8",
		x"77C377C277C177C0FFFFFFFFFFFFFFFF77BF77BE77BD77BC77BB77BA77B977B8",
		x"77D377D277D177D077CF77CE77CD77CC77CB77CA77C977C877C777C677C577C4",
		x"77E377E277E177E077DF77DE77DD77DC77DB77DA77D977D877D777D677D577D4",
		x"77F377F277F177F077EF77EE77ED77EC77EB77EA77E977E877E777E677E577E4",
		x"FFFFFFFFFFFFFFFF77FF77FE77FD77FC77FB77FA77F977F877F777F677F577F4",
		x"780F780E780D780C780B780A7809780878077806780578047803780278017800",
		x"781F781E781D781C781B781A7819781878177816781578147813781278117810",
		x"782F782E782D782C782B782A7829782878277826782578247823782278217820",
		x"783F783E783D783C783B783A7839783878377836783578347833783278317830",
		x"784B784A7849784878477846784578447843784278417840FFFFFFFFFFFFFFFF",
		x"785B785A7859785878577856785578547853785278517850784F784E784D784C",
		x"786B786A7869786878677866786578647863786278617860785F785E785D785C",
		x"787B787A7879787878777876787578747873787278717870786F786E786D786C",
		x"78877886788578847883788278817880FFFFFFFFFFFFFFFF787F787E787D787C",
		x"78977896789578947893789278917890788F788E788D788C788B788A78897888",
		x"78A778A678A578A478A378A278A178A0789F789E789D789C789B789A78997898",
		x"78B778B678B578B478B378B278B178B078AF78AE78AD78AC78AB78AA78A978A8",
		x"78C378C278C178C0FFFFFFFFFFFFFFFF78BF78BE78BD78BC78BB78BA78B978B8",
		x"78D378D278D178D078CF78CE78CD78CC78CB78CA78C978C878C778C678C578C4",
		x"78E378E278E178E078DF78DE78DD78DC78DB78DA78D978D878D778D678D578D4",
		x"78F378F278F178F078EF78EE78ED78EC78EB78EA78E978E878E778E678E578E4",
		x"FFFFFFFFFFFFFFFF78FF78FE78FD78FC78FB78FA78F978F878F778F678F578F4",
		x"790F790E790D790C790B790A7909790879077906790579047903790279017900",
		x"791F791E791D791C791B791A7919791879177916791579147913791279117910",
		x"792F792E792D792C792B792A7929792879277926792579247923792279217920",
		x"793F793E793D793C793B793A7939793879377936793579347933793279317930",
		x"794B794A7949794879477946794579447943794279417940FFFFFFFFFFFFFFFF",
		x"795B795A7959795879577956795579547953795279517950794F794E794D794C",
		x"796B796A7969796879677966796579647963796279617960795F795E795D795C",
		x"797B797A7979797879777976797579747973797279717970796F796E796D796C",
		x"79877986798579847983798279817980FFFFFFFFFFFFFFFF797F797E797D797C",
		x"79977996799579947993799279917990798F798E798D798C798B798A79897988",
		x"79A779A679A579A479A379A279A179A0799F799E799D799C799B799A79997998",
		x"79B779B679B579B479B379B279B179B079AF79AE79AD79AC79AB79AA79A979A8",
		x"79C379C279C179C0FFFFFFFFFFFFFFFF79BF79BE79BD79BC79BB79BA79B979B8",
		x"79D379D279D179D079CF79CE79CD79CC79CB79CA79C979C879C779C679C579C4",
		x"79E379E279E179E079DF79DE79DD79DC79DB79DA79D979D879D779D679D579D4",
		x"79F379F279F179F079EF79EE79ED79EC79EB79EA79E979E879E779E679E579E4",
		x"FFFFFFFFFFFFFFFF79FF79FE79FD79FC79FB79FA79F979F879F779F679F579F4",
		x"7A0F7A0E7A0D7A0C7A0B7A0A7A097A087A077A067A057A047A037A027A017A00",
		x"7A1F7A1E7A1D7A1C7A1B7A1A7A197A187A177A167A157A147A137A127A117A10",
		x"7A2F7A2E7A2D7A2C7A2B7A2A7A297A287A277A267A257A247A237A227A217A20",
		x"7A3F7A3E7A3D7A3C7A3B7A3A7A397A387A377A367A357A347A337A327A317A30",
		x"7A4B7A4A7A497A487A477A467A457A447A437A427A417A40FFFFFFFFFFFFFFFF",
		x"7A5B7A5A7A597A587A577A567A557A547A537A527A517A507A4F7A4E7A4D7A4C",
		x"7A6B7A6A7A697A687A677A667A657A647A637A627A617A607A5F7A5E7A5D7A5C",
		x"7A7B7A7A7A797A787A777A767A757A747A737A727A717A707A6F7A6E7A6D7A6C",
		x"7A877A867A857A847A837A827A817A80FFFFFFFFFFFFFFFF7A7F7A7E7A7D7A7C",
		x"7A977A967A957A947A937A927A917A907A8F7A8E7A8D7A8C7A8B7A8A7A897A88",
		x"7AA77AA67AA57AA47AA37AA27AA17AA07A9F7A9E7A9D7A9C7A9B7A9A7A997A98",
		x"7AB77AB67AB57AB47AB37AB27AB17AB07AAF7AAE7AAD7AAC7AAB7AAA7AA97AA8",
		x"7AC37AC27AC17AC0FFFFFFFFFFFFFFFF7ABF7ABE7ABD7ABC7ABB7ABA7AB97AB8",
		x"7AD37AD27AD17AD07ACF7ACE7ACD7ACC7ACB7ACA7AC97AC87AC77AC67AC57AC4",
		x"7AE37AE27AE17AE07ADF7ADE7ADD7ADC7ADB7ADA7AD97AD87AD77AD67AD57AD4",
		x"7AF37AF27AF17AF07AEF7AEE7AED7AEC7AEB7AEA7AE97AE87AE77AE67AE57AE4",
		x"FFFFFFFFFFFFFFFF7AFF7AFE7AFD7AFC7AFB7AFA7AF97AF87AF77AF67AF57AF4",
		x"7B0F7B0E7B0D7B0C7B0B7B0A7B097B087B077B067B057B047B037B027B017B00",
		x"7B1F7B1E7B1D7B1C7B1B7B1A7B197B187B177B167B157B147B137B127B117B10",
		x"7B2F7B2E7B2D7B2C7B2B7B2A7B297B287B277B267B257B247B237B227B217B20",
		x"7B3F7B3E7B3D7B3C7B3B7B3A7B397B387B377B367B357B347B337B327B317B30",
		x"7B4B7B4A7B497B487B477B467B457B447B437B427B417B40FFFFFFFFFFFFFFFF",
		x"7B5B7B5A7B597B587B577B567B557B547B537B527B517B507B4F7B4E7B4D7B4C",
		x"7B6B7B6A7B697B687B677B667B657B647B637B627B617B607B5F7B5E7B5D7B5C",
		x"7B7B7B7A7B797B787B777B767B757B747B737B727B717B707B6F7B6E7B6D7B6C",
		x"7B877B867B857B847B837B827B817B80FFFFFFFFFFFFFFFF7B7F7B7E7B7D7B7C",
		x"7B977B967B957B947B937B927B917B907B8F7B8E7B8D7B8C7B8B7B8A7B897B88",
		x"7BA77BA67BA57BA47BA37BA27BA17BA07B9F7B9E7B9D7B9C7B9B7B9A7B997B98",
		x"7BB77BB67BB57BB47BB37BB27BB17BB07BAF7BAE7BAD7BAC7BAB7BAA7BA97BA8",
		x"7BC37BC27BC17BC0FFFFFFFFFFFFFFFF7BBF7BBE7BBD7BBC7BBB7BBA7BB97BB8",
		x"7BD37BD27BD17BD07BCF7BCE7BCD7BCC7BCB7BCA7BC97BC87BC77BC67BC57BC4",
		x"7BE37BE27BE17BE07BDF7BDE7BDD7BDC7BDB7BDA7BD97BD87BD77BD67BD57BD4",
		x"7BF37BF27BF17BF07BEF7BEE7BED7BEC7BEB7BEA7BE97BE87BE77BE67BE57BE4",
		x"FFFFFFFFFFFFFFFF7BFF7BFE7BFD7BFC7BFB7BFA7BF97BF87BF77BF67BF57BF4",
		x"7C0F7C0E7C0D7C0C7C0B7C0A7C097C087C077C067C057C047C037C027C017C00",
		x"7C1F7C1E7C1D7C1C7C1B7C1A7C197C187C177C167C157C147C137C127C117C10",
		x"7C2F7C2E7C2D7C2C7C2B7C2A7C297C287C277C267C257C247C237C227C217C20",
		x"7C3F7C3E7C3D7C3C7C3B7C3A7C397C387C377C367C357C347C337C327C317C30",
		x"7C4B7C4A7C497C487C477C467C457C447C437C427C417C40FFFFFFFFFFFFFFFF",
		x"7C5B7C5A7C597C587C577C567C557C547C537C527C517C507C4F7C4E7C4D7C4C",
		x"7C6B7C6A7C697C687C677C667C657C647C637C627C617C607C5F7C5E7C5D7C5C",
		x"7C7B7C7A7C797C787C777C767C757C747C737C727C717C707C6F7C6E7C6D7C6C",
		x"7C877C867C857C847C837C827C817C80FFFFFFFFFFFFFFFF7C7F7C7E7C7D7C7C",
		x"7C977C967C957C947C937C927C917C907C8F7C8E7C8D7C8C7C8B7C8A7C897C88",
		x"7CA77CA67CA57CA47CA37CA27CA17CA07C9F7C9E7C9D7C9C7C9B7C9A7C997C98",
		x"7CB77CB67CB57CB47CB37CB27CB17CB07CAF7CAE7CAD7CAC7CAB7CAA7CA97CA8",
		x"7CC37CC27CC17CC0FFFFFFFFFFFFFFFF7CBF7CBE7CBD7CBC7CBB7CBA7CB97CB8",
		x"7CD37CD27CD17CD07CCF7CCE7CCD7CCC7CCB7CCA7CC97CC87CC77CC67CC57CC4",
		x"7CE37CE27CE17CE07CDF7CDE7CDD7CDC7CDB7CDA7CD97CD87CD77CD67CD57CD4",
		x"7CF37CF27CF17CF07CEF7CEE7CED7CEC7CEB7CEA7CE97CE87CE77CE67CE57CE4",
		x"FFFFFFFFFFFFFFFF7CFF7CFE7CFD7CFC7CFB7CFA7CF97CF87CF77CF67CF57CF4",
		x"7D0F7D0E7D0D7D0C7D0B7D0A7D097D087D077D067D057D047D037D027D017D00",
		x"7D1F7D1E7D1D7D1C7D1B7D1A7D197D187D177D167D157D147D137D127D117D10",
		x"7D2F7D2E7D2D7D2C7D2B7D2A7D297D287D277D267D257D247D237D227D217D20",
		x"7D3F7D3E7D3D7D3C7D3B7D3A7D397D387D377D367D357D347D337D327D317D30",
		x"7D4B7D4A7D497D487D477D467D457D447D437D427D417D40FFFFFFFFFFFFFFFF",
		x"7D5B7D5A7D597D587D577D567D557D547D537D527D517D507D4F7D4E7D4D7D4C",
		x"7D6B7D6A7D697D687D677D667D657D647D637D627D617D607D5F7D5E7D5D7D5C",
		x"7D7B7D7A7D797D787D777D767D757D747D737D727D717D707D6F7D6E7D6D7D6C",
		x"7D877D867D857D847D837D827D817D80FFFFFFFFFFFFFFFF7D7F7D7E7D7D7D7C",
		x"7D977D967D957D947D937D927D917D907D8F7D8E7D8D7D8C7D8B7D8A7D897D88",
		x"7DA77DA67DA57DA47DA37DA27DA17DA07D9F7D9E7D9D7D9C7D9B7D9A7D997D98",
		x"7DB77DB67DB57DB47DB37DB27DB17DB07DAF7DAE7DAD7DAC7DAB7DAA7DA97DA8",
		x"7DC37DC27DC17DC0FFFFFFFFFFFFFFFF7DBF7DBE7DBD7DBC7DBB7DBA7DB97DB8",
		x"7DD37DD27DD17DD07DCF7DCE7DCD7DCC7DCB7DCA7DC97DC87DC77DC67DC57DC4",
		x"7DE37DE27DE17DE07DDF7DDE7DDD7DDC7DDB7DDA7DD97DD87DD77DD67DD57DD4",
		x"7DF37DF27DF17DF07DEF7DEE7DED7DEC7DEB7DEA7DE97DE87DE77DE67DE57DE4",
		x"FFFFFFFFFFFFFFFF7DFF7DFE7DFD7DFC7DFB7DFA7DF97DF87DF77DF67DF57DF4",
		x"7E0F7E0E7E0D7E0C7E0B7E0A7E097E087E077E067E057E047E037E027E017E00",
		x"7E1F7E1E7E1D7E1C7E1B7E1A7E197E187E177E167E157E147E137E127E117E10",
		x"7E2F7E2E7E2D7E2C7E2B7E2A7E297E287E277E267E257E247E237E227E217E20",
		x"7E3F7E3E7E3D7E3C7E3B7E3A7E397E387E377E367E357E347E337E327E317E30",
		x"7E4B7E4A7E497E487E477E467E457E447E437E427E417E40FFFFFFFFFFFFFFFF",
		x"7E5B7E5A7E597E587E577E567E557E547E537E527E517E507E4F7E4E7E4D7E4C",
		x"7E6B7E6A7E697E687E677E667E657E647E637E627E617E607E5F7E5E7E5D7E5C",
		x"7E7B7E7A7E797E787E777E767E757E747E737E727E717E707E6F7E6E7E6D7E6C",
		x"7E877E867E857E847E837E827E817E80FFFFFFFFFFFFFFFF7E7F7E7E7E7D7E7C",
		x"7E977E967E957E947E937E927E917E907E8F7E8E7E8D7E8C7E8B7E8A7E897E88",
		x"7EA77EA67EA57EA47EA37EA27EA17EA07E9F7E9E7E9D7E9C7E9B7E9A7E997E98",
		x"7EB77EB67EB57EB47EB37EB27EB17EB07EAF7EAE7EAD7EAC7EAB7EAA7EA97EA8",
		x"7EC37EC27EC17EC0FFFFFFFFFFFFFFFF7EBF7EBE7EBD7EBC7EBB7EBA7EB97EB8",
		x"7ED37ED27ED17ED07ECF7ECE7ECD7ECC7ECB7ECA7EC97EC87EC77EC67EC57EC4",
		x"7EE37EE27EE17EE07EDF7EDE7EDD7EDC7EDB7EDA7ED97ED87ED77ED67ED57ED4",
		x"7EF37EF27EF17EF07EEF7EEE7EED7EEC7EEB7EEA7EE97EE87EE77EE67EE57EE4",
		x"FFFFFFFFFFFFFFFF7EFF7EFE7EFD7EFC7EFB7EFA7EF97EF87EF77EF67EF57EF4",
		x"7F0F7F0E7F0D7F0C7F0B7F0A7F097F087F077F067F057F047F037F027F017F00",
		x"7F1F7F1E7F1D7F1C7F1B7F1A7F197F187F177F167F157F147F137F127F117F10",
		x"7F2F7F2E7F2D7F2C7F2B7F2A7F297F287F277F267F257F247F237F227F217F20",
		x"7F3F7F3E7F3D7F3C7F3B7F3A7F397F387F377F367F357F347F337F327F317F30",
		x"7F4B7F4A7F497F487F477F467F457F447F437F427F417F40FFFFFFFFFFFFFFFF",
		x"7F5B7F5A7F597F587F577F567F557F547F537F527F517F507F4F7F4E7F4D7F4C",
		x"7F6B7F6A7F697F687F677F667F657F647F637F627F617F607F5F7F5E7F5D7F5C",
		x"7F7B7F7A7F797F787F777F767F757F747F737F727F717F707F6F7F6E7F6D7F6C",
		x"7F877F867F857F847F837F827F817F80FFFFFFFFFFFFFFFF7F7F7F7E7F7D7F7C",
		x"7F977F967F957F947F937F927F917F907F8F7F8E7F8D7F8C7F8B7F8A7F897F88",
		x"7FA77FA67FA57FA47FA37FA27FA17FA07F9F7F9E7F9D7F9C7F9B7F9A7F997F98",
		x"7FB77FB67FB57FB47FB37FB27FB17FB07FAF7FAE7FAD7FAC7FAB7FAA7FA97FA8",
		x"7FC37FC27FC17FC0FFFFFFFFFFFFFFFF7FBF7FBE7FBD7FBC7FBB7FBA7FB97FB8",
		x"7FD37FD27FD17FD07FCF7FCE7FCD7FCC7FCB7FCA7FC97FC87FC77FC67FC57FC4",
		x"7FE37FE27FE17FE07FDF7FDE7FDD7FDC7FDB7FDA7FD97FD87FD77FD67FD57FD4",
		x"7FF37FF27FF17FF07FEF7FEE7FED7FEC7FEB7FEA7FE97FE87FE77FE67FE57FE4",
		x"FFFFFFFFFFFFFFFF7FFF7FFE7FFD7FFC7FFB7FFA7FF97FF87FF77FF67FF57FF4",
		x"800F800E800D800C800B800A8009800880078006800580048003800280018000",
		x"801F801E801D801C801B801A8019801880178016801580148013801280118010",
		x"802F802E802D802C802B802A8029802880278026802580248023802280218020",
		x"803F803E803D803C803B803A8039803880378036803580348033803280318030",
		x"804B804A8049804880478046804580448043804280418040FFFFFFFFFFFFFFFF",
		x"805B805A8059805880578056805580548053805280518050804F804E804D804C",
		x"806B806A8069806880678066806580648063806280618060805F805E805D805C",
		x"807B807A8079807880778076807580748073807280718070806F806E806D806C",
		x"80878086808580848083808280818080FFFFFFFFFFFFFFFF807F807E807D807C",
		x"80978096809580948093809280918090808F808E808D808C808B808A80898088",
		x"80A780A680A580A480A380A280A180A0809F809E809D809C809B809A80998098",
		x"80B780B680B580B480B380B280B180B080AF80AE80AD80AC80AB80AA80A980A8",
		x"80C380C280C180C0FFFFFFFFFFFFFFFF80BF80BE80BD80BC80BB80BA80B980B8",
		x"80D380D280D180D080CF80CE80CD80CC80CB80CA80C980C880C780C680C580C4",
		x"80E380E280E180E080DF80DE80DD80DC80DB80DA80D980D880D780D680D580D4",
		x"80F380F280F180F080EF80EE80ED80EC80EB80EA80E980E880E780E680E580E4",
		x"FFFFFFFFFFFFFFFF80FF80FE80FD80FC80FB80FA80F980F880F780F680F580F4",
		x"810F810E810D810C810B810A8109810881078106810581048103810281018100",
		x"811F811E811D811C811B811A8119811881178116811581148113811281118110",
		x"812F812E812D812C812B812A8129812881278126812581248123812281218120",
		x"813F813E813D813C813B813A8139813881378136813581348133813281318130",
		x"814B814A8149814881478146814581448143814281418140FFFFFFFFFFFFFFFF",
		x"815B815A8159815881578156815581548153815281518150814F814E814D814C",
		x"816B816A8169816881678166816581648163816281618160815F815E815D815C",
		x"817B817A8179817881778176817581748173817281718170816F816E816D816C",
		x"81878186818581848183818281818180FFFFFFFFFFFFFFFF817F817E817D817C",
		x"81978196819581948193819281918190818F818E818D818C818B818A81898188",
		x"81A781A681A581A481A381A281A181A0819F819E819D819C819B819A81998198",
		x"81B781B681B581B481B381B281B181B081AF81AE81AD81AC81AB81AA81A981A8",
		x"81C381C281C181C0FFFFFFFFFFFFFFFF81BF81BE81BD81BC81BB81BA81B981B8",
		x"81D381D281D181D081CF81CE81CD81CC81CB81CA81C981C881C781C681C581C4",
		x"81E381E281E181E081DF81DE81DD81DC81DB81DA81D981D881D781D681D581D4",
		x"81F381F281F181F081EF81EE81ED81EC81EB81EA81E981E881E781E681E581E4",
		x"FFFFFFFFFFFFFFFF81FF81FE81FD81FC81FB81FA81F981F881F781F681F581F4",
		x"820F820E820D820C820B820A8209820882078206820582048203820282018200",
		x"821F821E821D821C821B821A8219821882178216821582148213821282118210",
		x"822F822E822D822C822B822A8229822882278226822582248223822282218220",
		x"823F823E823D823C823B823A8239823882378236823582348233823282318230",
		x"824B824A8249824882478246824582448243824282418240FFFFFFFFFFFFFFFF",
		x"825B825A8259825882578256825582548253825282518250824F824E824D824C",
		x"826B826A8269826882678266826582648263826282618260825F825E825D825C",
		x"827B827A8279827882778276827582748273827282718270826F826E826D826C",
		x"82878286828582848283828282818280FFFFFFFFFFFFFFFF827F827E827D827C",
		x"82978296829582948293829282918290828F828E828D828C828B828A82898288",
		x"82A782A682A582A482A382A282A182A0829F829E829D829C829B829A82998298",
		x"82B782B682B582B482B382B282B182B082AF82AE82AD82AC82AB82AA82A982A8",
		x"82C382C282C182C0FFFFFFFFFFFFFFFF82BF82BE82BD82BC82BB82BA82B982B8",
		x"82D382D282D182D082CF82CE82CD82CC82CB82CA82C982C882C782C682C582C4",
		x"82E382E282E182E082DF82DE82DD82DC82DB82DA82D982D882D782D682D582D4",
		x"82F382F282F182F082EF82EE82ED82EC82EB82EA82E982E882E782E682E582E4",
		x"FFFFFFFFFFFFFFFF82FF82FE82FD82FC82FB82FA82F982F882F782F682F582F4",
		x"830F830E830D830C830B830A8309830883078306830583048303830283018300",
		x"831F831E831D831C831B831A8319831883178316831583148313831283118310",
		x"832F832E832D832C832B832A8329832883278326832583248323832283218320",
		x"833F833E833D833C833B833A8339833883378336833583348333833283318330",
		x"834B834A8349834883478346834583448343834283418340FFFFFFFFFFFFFFFF",
		x"835B835A8359835883578356835583548353835283518350834F834E834D834C",
		x"836B836A8369836883678366836583648363836283618360835F835E835D835C",
		x"837B837A8379837883778376837583748373837283718370836F836E836D836C",
		x"83878386838583848383838283818380FFFFFFFFFFFFFFFF837F837E837D837C",
		x"83978396839583948393839283918390838F838E838D838C838B838A83898388",
		x"83A783A683A583A483A383A283A183A0839F839E839D839C839B839A83998398",
		x"83B783B683B583B483B383B283B183B083AF83AE83AD83AC83AB83AA83A983A8",
		x"83C383C283C183C0FFFFFFFFFFFFFFFF83BF83BE83BD83BC83BB83BA83B983B8",
		x"83D383D283D183D083CF83CE83CD83CC83CB83CA83C983C883C783C683C583C4",
		x"83E383E283E183E083DF83DE83DD83DC83DB83DA83D983D883D783D683D583D4",
		x"83F383F283F183F083EF83EE83ED83EC83EB83EA83E983E883E783E683E583E4",
		x"FFFFFFFFFFFFFFFF83FF83FE83FD83FC83FB83FA83F983F883F783F683F583F4",
		x"840F840E840D840C840B840A8409840884078406840584048403840284018400",
		x"841F841E841D841C841B841A8419841884178416841584148413841284118410",
		x"842F842E842D842C842B842A8429842884278426842584248423842284218420",
		x"843F843E843D843C843B843A8439843884378436843584348433843284318430",
		x"844B844A8449844884478446844584448443844284418440FFFFFFFFFFFFFFFF",
		x"845B845A8459845884578456845584548453845284518450844F844E844D844C",
		x"846B846A8469846884678466846584648463846284618460845F845E845D845C",
		x"847B847A8479847884778476847584748473847284718470846F846E846D846C",
		x"84878486848584848483848284818480FFFFFFFFFFFFFFFF847F847E847D847C",
		x"84978496849584948493849284918490848F848E848D848C848B848A84898488",
		x"84A784A684A584A484A384A284A184A0849F849E849D849C849B849A84998498",
		x"84B784B684B584B484B384B284B184B084AF84AE84AD84AC84AB84AA84A984A8",
		x"84C384C284C184C0FFFFFFFFFFFFFFFF84BF84BE84BD84BC84BB84BA84B984B8",
		x"84D384D284D184D084CF84CE84CD84CC84CB84CA84C984C884C784C684C584C4",
		x"84E384E284E184E084DF84DE84DD84DC84DB84DA84D984D884D784D684D584D4",
		x"84F384F284F184F084EF84EE84ED84EC84EB84EA84E984E884E784E684E584E4",
		x"FFFFFFFFFFFFFFFF84FF84FE84FD84FC84FB84FA84F984F884F784F684F584F4",
		x"850F850E850D850C850B850A8509850885078506850585048503850285018500",
		x"851F851E851D851C851B851A8519851885178516851585148513851285118510",
		x"852F852E852D852C852B852A8529852885278526852585248523852285218520",
		x"853F853E853D853C853B853A8539853885378536853585348533853285318530",
		x"854B854A8549854885478546854585448543854285418540FFFFFFFFFFFFFFFF",
		x"855B855A8559855885578556855585548553855285518550854F854E854D854C",
		x"856B856A8569856885678566856585648563856285618560855F855E855D855C",
		x"857B857A8579857885778576857585748573857285718570856F856E856D856C",
		x"85878586858585848583858285818580FFFFFFFFFFFFFFFF857F857E857D857C",
		x"85978596859585948593859285918590858F858E858D858C858B858A85898588",
		x"85A785A685A585A485A385A285A185A0859F859E859D859C859B859A85998598",
		x"85B785B685B585B485B385B285B185B085AF85AE85AD85AC85AB85AA85A985A8",
		x"85C385C285C185C0FFFFFFFFFFFFFFFF85BF85BE85BD85BC85BB85BA85B985B8",
		x"85D385D285D185D085CF85CE85CD85CC85CB85CA85C985C885C785C685C585C4",
		x"85E385E285E185E085DF85DE85DD85DC85DB85DA85D985D885D785D685D585D4",
		x"85F385F285F185F085EF85EE85ED85EC85EB85EA85E985E885E785E685E585E4",
		x"FFFFFFFFFFFFFFFF85FF85FE85FD85FC85FB85FA85F985F885F785F685F585F4",
		x"860F860E860D860C860B860A8609860886078606860586048603860286018600",
		x"861F861E861D861C861B861A8619861886178616861586148613861286118610",
		x"862F862E862D862C862B862A8629862886278626862586248623862286218620",
		x"863F863E863D863C863B863A8639863886378636863586348633863286318630",
		x"864B864A8649864886478646864586448643864286418640FFFFFFFFFFFFFFFF",
		x"865B865A8659865886578656865586548653865286518650864F864E864D864C",
		x"866B866A8669866886678666866586648663866286618660865F865E865D865C",
		x"867B867A8679867886778676867586748673867286718670866F866E866D866C",
		x"86878686868586848683868286818680FFFFFFFFFFFFFFFF867F867E867D867C",
		x"86978696869586948693869286918690868F868E868D868C868B868A86898688",
		x"86A786A686A586A486A386A286A186A0869F869E869D869C869B869A86998698",
		x"86B786B686B586B486B386B286B186B086AF86AE86AD86AC86AB86AA86A986A8",
		x"86C386C286C186C0FFFFFFFFFFFFFFFF86BF86BE86BD86BC86BB86BA86B986B8",
		x"86D386D286D186D086CF86CE86CD86CC86CB86CA86C986C886C786C686C586C4",
		x"86E386E286E186E086DF86DE86DD86DC86DB86DA86D986D886D786D686D586D4",
		x"86F386F286F186F086EF86EE86ED86EC86EB86EA86E986E886E786E686E586E4",
		x"FFFFFFFFFFFFFFFF86FF86FE86FD86FC86FB86FA86F986F886F786F686F586F4",
		x"870F870E870D870C870B870A8709870887078706870587048703870287018700",
		x"871F871E871D871C871B871A8719871887178716871587148713871287118710",
		x"872F872E872D872C872B872A8729872887278726872587248723872287218720",
		x"873F873E873D873C873B873A8739873887378736873587348733873287318730",
		x"874B874A8749874887478746874587448743874287418740FFFFFFFFFFFFFFFF",
		x"875B875A8759875887578756875587548753875287518750874F874E874D874C",
		x"876B876A8769876887678766876587648763876287618760875F875E875D875C",
		x"877B877A8779877887778776877587748773877287718770876F876E876D876C",
		x"87878786878587848783878287818780FFFFFFFFFFFFFFFF877F877E877D877C",
		x"87978796879587948793879287918790878F878E878D878C878B878A87898788",
		x"87A787A687A587A487A387A287A187A0879F879E879D879C879B879A87998798",
		x"87B787B687B587B487B387B287B187B087AF87AE87AD87AC87AB87AA87A987A8",
		x"87C387C287C187C0FFFFFFFFFFFFFFFF87BF87BE87BD87BC87BB87BA87B987B8",
		x"87D387D287D187D087CF87CE87CD87CC87CB87CA87C987C887C787C687C587C4",
		x"87E387E287E187E087DF87DE87DD87DC87DB87DA87D987D887D787D687D587D4",
		x"87F387F287F187F087EF87EE87ED87EC87EB87EA87E987E887E787E687E587E4",
		x"FFFFFFFFFFFFFFFF87FF87FE87FD87FC87FB87FA87F987F887F787F687F587F4",
		x"880F880E880D880C880B880A8809880888078806880588048803880288018800",
		x"881F881E881D881C881B881A8819881888178816881588148813881288118810",
		x"882F882E882D882C882B882A8829882888278826882588248823882288218820",
		x"883F883E883D883C883B883A8839883888378836883588348833883288318830",
		x"884B884A8849884888478846884588448843884288418840FFFFFFFFFFFFFFFF",
		x"885B885A8859885888578856885588548853885288518850884F884E884D884C",
		x"886B886A8869886888678866886588648863886288618860885F885E885D885C",
		x"887B887A8879887888778876887588748873887288718870886F886E886D886C",
		x"88878886888588848883888288818880FFFFFFFFFFFFFFFF887F887E887D887C",
		x"88978896889588948893889288918890888F888E888D888C888B888A88898888",
		x"88A788A688A588A488A388A288A188A0889F889E889D889C889B889A88998898",
		x"88B788B688B588B488B388B288B188B088AF88AE88AD88AC88AB88AA88A988A8",
		x"88C388C288C188C0FFFFFFFFFFFFFFFF88BF88BE88BD88BC88BB88BA88B988B8",
		x"88D388D288D188D088CF88CE88CD88CC88CB88CA88C988C888C788C688C588C4",
		x"88E388E288E188E088DF88DE88DD88DC88DB88DA88D988D888D788D688D588D4",
		x"88F388F288F188F088EF88EE88ED88EC88EB88EA88E988E888E788E688E588E4",
		x"FFFFFFFFFFFFFFFF88FF88FE88FD88FC88FB88FA88F988F888F788F688F588F4",
		x"890F890E890D890C890B890A8909890889078906890589048903890289018900",
		x"891F891E891D891C891B891A8919891889178916891589148913891289118910",
		x"892F892E892D892C892B892A8929892889278926892589248923892289218920",
		x"893F893E893D893C893B893A8939893889378936893589348933893289318930",
		x"894B894A8949894889478946894589448943894289418940FFFFFFFFFFFFFFFF",
		x"895B895A8959895889578956895589548953895289518950894F894E894D894C",
		x"896B896A8969896889678966896589648963896289618960895F895E895D895C",
		x"897B897A8979897889778976897589748973897289718970896F896E896D896C",
		x"89878986898589848983898289818980FFFFFFFFFFFFFFFF897F897E897D897C",
		x"89978996899589948993899289918990898F898E898D898C898B898A89898988",
		x"89A789A689A589A489A389A289A189A0899F899E899D899C899B899A89998998",
		x"89B789B689B589B489B389B289B189B089AF89AE89AD89AC89AB89AA89A989A8",
		x"89C389C289C189C0FFFFFFFFFFFFFFFF89BF89BE89BD89BC89BB89BA89B989B8",
		x"89D389D289D189D089CF89CE89CD89CC89CB89CA89C989C889C789C689C589C4",
		x"89E389E289E189E089DF89DE89DD89DC89DB89DA89D989D889D789D689D589D4",
		x"89F389F289F189F089EF89EE89ED89EC89EB89EA89E989E889E789E689E589E4",
		x"FFFFFFFFFFFFFFFF89FF89FE89FD89FC89FB89FA89F989F889F789F689F589F4",
		x"8A0F8A0E8A0D8A0C8A0B8A0A8A098A088A078A068A058A048A038A028A018A00",
		x"8A1F8A1E8A1D8A1C8A1B8A1A8A198A188A178A168A158A148A138A128A118A10",
		x"8A2F8A2E8A2D8A2C8A2B8A2A8A298A288A278A268A258A248A238A228A218A20",
		x"8A3F8A3E8A3D8A3C8A3B8A3A8A398A388A378A368A358A348A338A328A318A30",
		x"8A4B8A4A8A498A488A478A468A458A448A438A428A418A40FFFFFFFFFFFFFFFF",
		x"8A5B8A5A8A598A588A578A568A558A548A538A528A518A508A4F8A4E8A4D8A4C",
		x"8A6B8A6A8A698A688A678A668A658A648A638A628A618A608A5F8A5E8A5D8A5C",
		x"8A7B8A7A8A798A788A778A768A758A748A738A728A718A708A6F8A6E8A6D8A6C",
		x"8A878A868A858A848A838A828A818A80FFFFFFFFFFFFFFFF8A7F8A7E8A7D8A7C",
		x"8A978A968A958A948A938A928A918A908A8F8A8E8A8D8A8C8A8B8A8A8A898A88",
		x"8AA78AA68AA58AA48AA38AA28AA18AA08A9F8A9E8A9D8A9C8A9B8A9A8A998A98",
		x"8AB78AB68AB58AB48AB38AB28AB18AB08AAF8AAE8AAD8AAC8AAB8AAA8AA98AA8",
		x"8AC38AC28AC18AC0FFFFFFFFFFFFFFFF8ABF8ABE8ABD8ABC8ABB8ABA8AB98AB8",
		x"8AD38AD28AD18AD08ACF8ACE8ACD8ACC8ACB8ACA8AC98AC88AC78AC68AC58AC4",
		x"8AE38AE28AE18AE08ADF8ADE8ADD8ADC8ADB8ADA8AD98AD88AD78AD68AD58AD4",
		x"8AF38AF28AF18AF08AEF8AEE8AED8AEC8AEB8AEA8AE98AE88AE78AE68AE58AE4",
		x"FFFFFFFFFFFFFFFF8AFF8AFE8AFD8AFC8AFB8AFA8AF98AF88AF78AF68AF58AF4",
		x"8B0F8B0E8B0D8B0C8B0B8B0A8B098B088B078B068B058B048B038B028B018B00",
		x"8B1F8B1E8B1D8B1C8B1B8B1A8B198B188B178B168B158B148B138B128B118B10",
		x"8B2F8B2E8B2D8B2C8B2B8B2A8B298B288B278B268B258B248B238B228B218B20",
		x"8B3F8B3E8B3D8B3C8B3B8B3A8B398B388B378B368B358B348B338B328B318B30",
		x"8B4B8B4A8B498B488B478B468B458B448B438B428B418B40FFFFFFFFFFFFFFFF",
		x"8B5B8B5A8B598B588B578B568B558B548B538B528B518B508B4F8B4E8B4D8B4C",
		x"8B6B8B6A8B698B688B678B668B658B648B638B628B618B608B5F8B5E8B5D8B5C",
		x"8B7B8B7A8B798B788B778B768B758B748B738B728B718B708B6F8B6E8B6D8B6C",
		x"8B878B868B858B848B838B828B818B80FFFFFFFFFFFFFFFF8B7F8B7E8B7D8B7C",
		x"8B978B968B958B948B938B928B918B908B8F8B8E8B8D8B8C8B8B8B8A8B898B88",
		x"8BA78BA68BA58BA48BA38BA28BA18BA08B9F8B9E8B9D8B9C8B9B8B9A8B998B98",
		x"8BB78BB68BB58BB48BB38BB28BB18BB08BAF8BAE8BAD8BAC8BAB8BAA8BA98BA8",
		x"8BC38BC28BC18BC0FFFFFFFFFFFFFFFF8BBF8BBE8BBD8BBC8BBB8BBA8BB98BB8",
		x"8BD38BD28BD18BD08BCF8BCE8BCD8BCC8BCB8BCA8BC98BC88BC78BC68BC58BC4",
		x"8BE38BE28BE18BE08BDF8BDE8BDD8BDC8BDB8BDA8BD98BD88BD78BD68BD58BD4",
		x"8BF38BF28BF18BF08BEF8BEE8BED8BEC8BEB8BEA8BE98BE88BE78BE68BE58BE4",
		x"FFFFFFFFFFFFFFFF8BFF8BFE8BFD8BFC8BFB8BFA8BF98BF88BF78BF68BF58BF4",
		x"8C0F8C0E8C0D8C0C8C0B8C0A8C098C088C078C068C058C048C038C028C018C00",
		x"8C1F8C1E8C1D8C1C8C1B8C1A8C198C188C178C168C158C148C138C128C118C10",
		x"8C2F8C2E8C2D8C2C8C2B8C2A8C298C288C278C268C258C248C238C228C218C20",
		x"8C3F8C3E8C3D8C3C8C3B8C3A8C398C388C378C368C358C348C338C328C318C30",
		x"8C4B8C4A8C498C488C478C468C458C448C438C428C418C40FFFFFFFFFFFFFFFF",
		x"8C5B8C5A8C598C588C578C568C558C548C538C528C518C508C4F8C4E8C4D8C4C",
		x"8C6B8C6A8C698C688C678C668C658C648C638C628C618C608C5F8C5E8C5D8C5C",
		x"8C7B8C7A8C798C788C778C768C758C748C738C728C718C708C6F8C6E8C6D8C6C",
		x"8C878C868C858C848C838C828C818C80FFFFFFFFFFFFFFFF8C7F8C7E8C7D8C7C",
		x"8C978C968C958C948C938C928C918C908C8F8C8E8C8D8C8C8C8B8C8A8C898C88",
		x"8CA78CA68CA58CA48CA38CA28CA18CA08C9F8C9E8C9D8C9C8C9B8C9A8C998C98",
		x"8CB78CB68CB58CB48CB38CB28CB18CB08CAF8CAE8CAD8CAC8CAB8CAA8CA98CA8",
		x"8CC38CC28CC18CC0FFFFFFFFFFFFFFFF8CBF8CBE8CBD8CBC8CBB8CBA8CB98CB8",
		x"8CD38CD28CD18CD08CCF8CCE8CCD8CCC8CCB8CCA8CC98CC88CC78CC68CC58CC4",
		x"8CE38CE28CE18CE08CDF8CDE8CDD8CDC8CDB8CDA8CD98CD88CD78CD68CD58CD4",
		x"8CF38CF28CF18CF08CEF8CEE8CED8CEC8CEB8CEA8CE98CE88CE78CE68CE58CE4",
		x"FFFFFFFFFFFFFFFF8CFF8CFE8CFD8CFC8CFB8CFA8CF98CF88CF78CF68CF58CF4",
		x"8D0F8D0E8D0D8D0C8D0B8D0A8D098D088D078D068D058D048D038D028D018D00",
		x"8D1F8D1E8D1D8D1C8D1B8D1A8D198D188D178D168D158D148D138D128D118D10",
		x"8D2F8D2E8D2D8D2C8D2B8D2A8D298D288D278D268D258D248D238D228D218D20",
		x"8D3F8D3E8D3D8D3C8D3B8D3A8D398D388D378D368D358D348D338D328D318D30",
		x"8D4B8D4A8D498D488D478D468D458D448D438D428D418D40FFFFFFFFFFFFFFFF",
		x"8D5B8D5A8D598D588D578D568D558D548D538D528D518D508D4F8D4E8D4D8D4C",
		x"8D6B8D6A8D698D688D678D668D658D648D638D628D618D608D5F8D5E8D5D8D5C",
		x"8D7B8D7A8D798D788D778D768D758D748D738D728D718D708D6F8D6E8D6D8D6C",
		x"8D878D868D858D848D838D828D818D80FFFFFFFFFFFFFFFF8D7F8D7E8D7D8D7C",
		x"8D978D968D958D948D938D928D918D908D8F8D8E8D8D8D8C8D8B8D8A8D898D88",
		x"8DA78DA68DA58DA48DA38DA28DA18DA08D9F8D9E8D9D8D9C8D9B8D9A8D998D98",
		x"8DB78DB68DB58DB48DB38DB28DB18DB08DAF8DAE8DAD8DAC8DAB8DAA8DA98DA8",
		x"8DC38DC28DC18DC0FFFFFFFFFFFFFFFF8DBF8DBE8DBD8DBC8DBB8DBA8DB98DB8",
		x"8DD38DD28DD18DD08DCF8DCE8DCD8DCC8DCB8DCA8DC98DC88DC78DC68DC58DC4",
		x"8DE38DE28DE18DE08DDF8DDE8DDD8DDC8DDB8DDA8DD98DD88DD78DD68DD58DD4",
		x"8DF38DF28DF18DF08DEF8DEE8DED8DEC8DEB8DEA8DE98DE88DE78DE68DE58DE4",
		x"FFFFFFFFFFFFFFFF8DFF8DFE8DFD8DFC8DFB8DFA8DF98DF88DF78DF68DF58DF4",
		x"8E0F8E0E8E0D8E0C8E0B8E0A8E098E088E078E068E058E048E038E028E018E00",
		x"8E1F8E1E8E1D8E1C8E1B8E1A8E198E188E178E168E158E148E138E128E118E10",
		x"8E2F8E2E8E2D8E2C8E2B8E2A8E298E288E278E268E258E248E238E228E218E20",
		x"8E3F8E3E8E3D8E3C8E3B8E3A8E398E388E378E368E358E348E338E328E318E30",
		x"8E4B8E4A8E498E488E478E468E458E448E438E428E418E40FFFFFFFFFFFFFFFF",
		x"8E5B8E5A8E598E588E578E568E558E548E538E528E518E508E4F8E4E8E4D8E4C",
		x"8E6B8E6A8E698E688E678E668E658E648E638E628E618E608E5F8E5E8E5D8E5C",
		x"8E7B8E7A8E798E788E778E768E758E748E738E728E718E708E6F8E6E8E6D8E6C",
		x"8E878E868E858E848E838E828E818E80FFFFFFFFFFFFFFFF8E7F8E7E8E7D8E7C",
		x"8E978E968E958E948E938E928E918E908E8F8E8E8E8D8E8C8E8B8E8A8E898E88",
		x"8EA78EA68EA58EA48EA38EA28EA18EA08E9F8E9E8E9D8E9C8E9B8E9A8E998E98",
		x"8EB78EB68EB58EB48EB38EB28EB18EB08EAF8EAE8EAD8EAC8EAB8EAA8EA98EA8",
		x"8EC38EC28EC18EC0FFFFFFFFFFFFFFFF8EBF8EBE8EBD8EBC8EBB8EBA8EB98EB8",
		x"8ED38ED28ED18ED08ECF8ECE8ECD8ECC8ECB8ECA8EC98EC88EC78EC68EC58EC4",
		x"8EE38EE28EE18EE08EDF8EDE8EDD8EDC8EDB8EDA8ED98ED88ED78ED68ED58ED4",
		x"8EF38EF28EF18EF08EEF8EEE8EED8EEC8EEB8EEA8EE98EE88EE78EE68EE58EE4",
		x"FFFFFFFFFFFFFFFF8EFF8EFE8EFD8EFC8EFB8EFA8EF98EF88EF78EF68EF58EF4",
		x"8F0F8F0E8F0D8F0C8F0B8F0A8F098F088F078F068F058F048F038F028F018F00",
		x"8F1F8F1E8F1D8F1C8F1B8F1A8F198F188F178F168F158F148F138F128F118F10",
		x"8F2F8F2E8F2D8F2C8F2B8F2A8F298F288F278F268F258F248F238F228F218F20",
		x"8F3F8F3E8F3D8F3C8F3B8F3A8F398F388F378F368F358F348F338F328F318F30",
		x"8F4B8F4A8F498F488F478F468F458F448F438F428F418F40FFFFFFFFFFFFFFFF",
		x"8F5B8F5A8F598F588F578F568F558F548F538F528F518F508F4F8F4E8F4D8F4C",
		x"8F6B8F6A8F698F688F678F668F658F648F638F628F618F608F5F8F5E8F5D8F5C",
		x"8F7B8F7A8F798F788F778F768F758F748F738F728F718F708F6F8F6E8F6D8F6C",
		x"8F878F868F858F848F838F828F818F80FFFFFFFFFFFFFFFF8F7F8F7E8F7D8F7C",
		x"8F978F968F958F948F938F928F918F908F8F8F8E8F8D8F8C8F8B8F8A8F898F88",
		x"8FA78FA68FA58FA48FA38FA28FA18FA08F9F8F9E8F9D8F9C8F9B8F9A8F998F98",
		x"8FB78FB68FB58FB48FB38FB28FB18FB08FAF8FAE8FAD8FAC8FAB8FAA8FA98FA8",
		x"8FC38FC28FC18FC0FFFFFFFFFFFFFFFF8FBF8FBE8FBD8FBC8FBB8FBA8FB98FB8",
		x"8FD38FD28FD18FD08FCF8FCE8FCD8FCC8FCB8FCA8FC98FC88FC78FC68FC58FC4",
		x"8FE38FE28FE18FE08FDF8FDE8FDD8FDC8FDB8FDA8FD98FD88FD78FD68FD58FD4",
		x"8FF38FF28FF18FF08FEF8FEE8FED8FEC8FEB8FEA8FE98FE88FE78FE68FE58FE4",
		x"FFFFFFFFFFFFFFFF8FFF8FFE8FFD8FFC8FFB8FFA8FF98FF88FF78FF68FF58FF4",
		x"900F900E900D900C900B900A9009900890079006900590049003900290019000",
		x"901F901E901D901C901B901A9019901890179016901590149013901290119010",
		x"902F902E902D902C902B902A9029902890279026902590249023902290219020",
		x"903F903E903D903C903B903A9039903890379036903590349033903290319030",
		x"904B904A9049904890479046904590449043904290419040FFFFFFFFFFFFFFFF",
		x"905B905A9059905890579056905590549053905290519050904F904E904D904C",
		x"906B906A9069906890679066906590649063906290619060905F905E905D905C",
		x"907B907A9079907890779076907590749073907290719070906F906E906D906C",
		x"90879086908590849083908290819080FFFFFFFFFFFFFFFF907F907E907D907C",
		x"90979096909590949093909290919090908F908E908D908C908B908A90899088",
		x"90A790A690A590A490A390A290A190A0909F909E909D909C909B909A90999098",
		x"90B790B690B590B490B390B290B190B090AF90AE90AD90AC90AB90AA90A990A8",
		x"90C390C290C190C0FFFFFFFFFFFFFFFF90BF90BE90BD90BC90BB90BA90B990B8",
		x"90D390D290D190D090CF90CE90CD90CC90CB90CA90C990C890C790C690C590C4",
		x"90E390E290E190E090DF90DE90DD90DC90DB90DA90D990D890D790D690D590D4",
		x"90F390F290F190F090EF90EE90ED90EC90EB90EA90E990E890E790E690E590E4",
		x"FFFFFFFFFFFFFFFF90FF90FE90FD90FC90FB90FA90F990F890F790F690F590F4",
		x"910F910E910D910C910B910A9109910891079106910591049103910291019100",
		x"911F911E911D911C911B911A9119911891179116911591149113911291119110",
		x"912F912E912D912C912B912A9129912891279126912591249123912291219120",
		x"913F913E913D913C913B913A9139913891379136913591349133913291319130",
		x"914B914A9149914891479146914591449143914291419140FFFFFFFFFFFFFFFF",
		x"915B915A9159915891579156915591549153915291519150914F914E914D914C",
		x"916B916A9169916891679166916591649163916291619160915F915E915D915C",
		x"917B917A9179917891779176917591749173917291719170916F916E916D916C",
		x"91879186918591849183918291819180FFFFFFFFFFFFFFFF917F917E917D917C",
		x"91979196919591949193919291919190918F918E918D918C918B918A91899188",
		x"91A791A691A591A491A391A291A191A0919F919E919D919C919B919A91999198",
		x"91B791B691B591B491B391B291B191B091AF91AE91AD91AC91AB91AA91A991A8",
		x"91C391C291C191C0FFFFFFFFFFFFFFFF91BF91BE91BD91BC91BB91BA91B991B8",
		x"91D391D291D191D091CF91CE91CD91CC91CB91CA91C991C891C791C691C591C4",
		x"91E391E291E191E091DF91DE91DD91DC91DB91DA91D991D891D791D691D591D4",
		x"91F391F291F191F091EF91EE91ED91EC91EB91EA91E991E891E791E691E591E4",
		x"FFFFFFFFFFFFFFFF91FF91FE91FD91FC91FB91FA91F991F891F791F691F591F4",
		x"920F920E920D920C920B920A9209920892079206920592049203920292019200",
		x"921F921E921D921C921B921A9219921892179216921592149213921292119210",
		x"922F922E922D922C922B922A9229922892279226922592249223922292219220",
		x"923F923E923D923C923B923A9239923892379236923592349233923292319230",
		x"924B924A9249924892479246924592449243924292419240FFFFFFFFFFFFFFFF",
		x"925B925A9259925892579256925592549253925292519250924F924E924D924C",
		x"926B926A9269926892679266926592649263926292619260925F925E925D925C",
		x"927B927A9279927892779276927592749273927292719270926F926E926D926C",
		x"92879286928592849283928292819280FFFFFFFFFFFFFFFF927F927E927D927C",
		x"92979296929592949293929292919290928F928E928D928C928B928A92899288",
		x"92A792A692A592A492A392A292A192A0929F929E929D929C929B929A92999298",
		x"92B792B692B592B492B392B292B192B092AF92AE92AD92AC92AB92AA92A992A8",
		x"92C392C292C192C0FFFFFFFFFFFFFFFF92BF92BE92BD92BC92BB92BA92B992B8",
		x"92D392D292D192D092CF92CE92CD92CC92CB92CA92C992C892C792C692C592C4",
		x"92E392E292E192E092DF92DE92DD92DC92DB92DA92D992D892D792D692D592D4",
		x"92F392F292F192F092EF92EE92ED92EC92EB92EA92E992E892E792E692E592E4",
		x"FFFFFFFFFFFFFFFF92FF92FE92FD92FC92FB92FA92F992F892F792F692F592F4",
		x"930F930E930D930C930B930A9309930893079306930593049303930293019300",
		x"931F931E931D931C931B931A9319931893179316931593149313931293119310",
		x"932F932E932D932C932B932A9329932893279326932593249323932293219320",
		x"933F933E933D933C933B933A9339933893379336933593349333933293319330",
		x"934B934A9349934893479346934593449343934293419340FFFFFFFFFFFFFFFF",
		x"935B935A9359935893579356935593549353935293519350934F934E934D934C",
		x"936B936A9369936893679366936593649363936293619360935F935E935D935C",
		x"937B937A9379937893779376937593749373937293719370936F936E936D936C",
		x"93879386938593849383938293819380FFFFFFFFFFFFFFFF937F937E937D937C",
		x"93979396939593949393939293919390938F938E938D938C938B938A93899388",
		x"93A793A693A593A493A393A293A193A0939F939E939D939C939B939A93999398",
		x"93B793B693B593B493B393B293B193B093AF93AE93AD93AC93AB93AA93A993A8",
		x"93C393C293C193C0FFFFFFFFFFFFFFFF93BF93BE93BD93BC93BB93BA93B993B8",
		x"93D393D293D193D093CF93CE93CD93CC93CB93CA93C993C893C793C693C593C4",
		x"93E393E293E193E093DF93DE93DD93DC93DB93DA93D993D893D793D693D593D4",
		x"93F393F293F193F093EF93EE93ED93EC93EB93EA93E993E893E793E693E593E4",
		x"FFFFFFFFFFFFFFFF93FF93FE93FD93FC93FB93FA93F993F893F793F693F593F4",
		x"940F940E940D940C940B940A9409940894079406940594049403940294019400",
		x"941F941E941D941C941B941A9419941894179416941594149413941294119410",
		x"942F942E942D942C942B942A9429942894279426942594249423942294219420",
		x"943F943E943D943C943B943A9439943894379436943594349433943294319430",
		x"944B944A9449944894479446944594449443944294419440FFFFFFFFFFFFFFFF",
		x"945B945A9459945894579456945594549453945294519450944F944E944D944C",
		x"946B946A9469946894679466946594649463946294619460945F945E945D945C",
		x"947B947A9479947894779476947594749473947294719470946F946E946D946C",
		x"94879486948594849483948294819480FFFFFFFFFFFFFFFF947F947E947D947C",
		x"94979496949594949493949294919490948F948E948D948C948B948A94899488",
		x"94A794A694A594A494A394A294A194A0949F949E949D949C949B949A94999498",
		x"94B794B694B594B494B394B294B194B094AF94AE94AD94AC94AB94AA94A994A8",
		x"94C394C294C194C0FFFFFFFFFFFFFFFF94BF94BE94BD94BC94BB94BA94B994B8",
		x"94D394D294D194D094CF94CE94CD94CC94CB94CA94C994C894C794C694C594C4",
		x"94E394E294E194E094DF94DE94DD94DC94DB94DA94D994D894D794D694D594D4",
		x"94F394F294F194F094EF94EE94ED94EC94EB94EA94E994E894E794E694E594E4",
		x"FFFFFFFFFFFFFFFF94FF94FE94FD94FC94FB94FA94F994F894F794F694F594F4",
		x"950F950E950D950C950B950A9509950895079506950595049503950295019500",
		x"951F951E951D951C951B951A9519951895179516951595149513951295119510",
		x"952F952E952D952C952B952A9529952895279526952595249523952295219520",
		x"953F953E953D953C953B953A9539953895379536953595349533953295319530",
		x"954B954A9549954895479546954595449543954295419540FFFFFFFFFFFFFFFF",
		x"955B955A9559955895579556955595549553955295519550954F954E954D954C",
		x"956B956A9569956895679566956595649563956295619560955F955E955D955C",
		x"957B957A9579957895779576957595749573957295719570956F956E956D956C",
		x"95879586958595849583958295819580FFFFFFFFFFFFFFFF957F957E957D957C",
		x"95979596959595949593959295919590958F958E958D958C958B958A95899588",
		x"95A795A695A595A495A395A295A195A0959F959E959D959C959B959A95999598",
		x"95B795B695B595B495B395B295B195B095AF95AE95AD95AC95AB95AA95A995A8",
		x"95C395C295C195C0FFFFFFFFFFFFFFFF95BF95BE95BD95BC95BB95BA95B995B8",
		x"95D395D295D195D095CF95CE95CD95CC95CB95CA95C995C895C795C695C595C4",
		x"95E395E295E195E095DF95DE95DD95DC95DB95DA95D995D895D795D695D595D4",
		x"95F395F295F195F095EF95EE95ED95EC95EB95EA95E995E895E795E695E595E4",
		x"FFFFFFFFFFFFFFFF95FF95FE95FD95FC95FB95FA95F995F895F795F695F595F4",
		x"960F960E960D960C960B960A9609960896079606960596049603960296019600",
		x"961F961E961D961C961B961A9619961896179616961596149613961296119610",
		x"962F962E962D962C962B962A9629962896279626962596249623962296219620",
		x"963F963E963D963C963B963A9639963896379636963596349633963296319630",
		x"964B964A9649964896479646964596449643964296419640FFFFFFFFFFFFFFFF",
		x"965B965A9659965896579656965596549653965296519650964F964E964D964C",
		x"966B966A9669966896679666966596649663966296619660965F965E965D965C",
		x"967B967A9679967896779676967596749673967296719670966F966E966D966C",
		x"96879686968596849683968296819680FFFFFFFFFFFFFFFF967F967E967D967C",
		x"96979696969596949693969296919690968F968E968D968C968B968A96899688",
		x"96A796A696A596A496A396A296A196A0969F969E969D969C969B969A96999698",
		x"96B796B696B596B496B396B296B196B096AF96AE96AD96AC96AB96AA96A996A8",
		x"96C396C296C196C0FFFFFFFFFFFFFFFF96BF96BE96BD96BC96BB96BA96B996B8",
		x"96D396D296D196D096CF96CE96CD96CC96CB96CA96C996C896C796C696C596C4",
		x"96E396E296E196E096DF96DE96DD96DC96DB96DA96D996D896D796D696D596D4",
		x"96F396F296F196F096EF96EE96ED96EC96EB96EA96E996E896E796E696E596E4",
		x"FFFFFFFFFFFFFFFF96FF96FE96FD96FC96FB96FA96F996F896F796F696F596F4",
		x"970F970E970D970C970B970A9709970897079706970597049703970297019700",
		x"971F971E971D971C971B971A9719971897179716971597149713971297119710",
		x"972F972E972D972C972B972A9729972897279726972597249723972297219720",
		x"973F973E973D973C973B973A9739973897379736973597349733973297319730",
		x"974B974A9749974897479746974597449743974297419740FFFFFFFFFFFFFFFF",
		x"975B975A9759975897579756975597549753975297519750974F974E974D974C",
		x"976B976A9769976897679766976597649763976297619760975F975E975D975C",
		x"977B977A9779977897779776977597749773977297719770976F976E976D976C",
		x"97879786978597849783978297819780FFFFFFFFFFFFFFFF977F977E977D977C",
		x"97979796979597949793979297919790978F978E978D978C978B978A97899788",
		x"97A797A697A597A497A397A297A197A0979F979E979D979C979B979A97999798",
		x"97B797B697B597B497B397B297B197B097AF97AE97AD97AC97AB97AA97A997A8",
		x"97C397C297C197C0FFFFFFFFFFFFFFFF97BF97BE97BD97BC97BB97BA97B997B8",
		x"97D397D297D197D097CF97CE97CD97CC97CB97CA97C997C897C797C697C597C4",
		x"97E397E297E197E097DF97DE97DD97DC97DB97DA97D997D897D797D697D597D4",
		x"97F397F297F197F097EF97EE97ED97EC97EB97EA97E997E897E797E697E597E4",
		x"FFFFFFFFFFFFFFFF97FF97FE97FD97FC97FB97FA97F997F897F797F697F597F4",
		x"980F980E980D980C980B980A9809980898079806980598049803980298019800",
		x"981F981E981D981C981B981A9819981898179816981598149813981298119810",
		x"982F982E982D982C982B982A9829982898279826982598249823982298219820",
		x"983F983E983D983C983B983A9839983898379836983598349833983298319830",
		x"984B984A9849984898479846984598449843984298419840FFFFFFFFFFFFFFFF",
		x"985B985A9859985898579856985598549853985298519850984F984E984D984C",
		x"986B986A9869986898679866986598649863986298619860985F985E985D985C",
		x"987B987A9879987898779876987598749873987298719870986F986E986D986C",
		x"98879886988598849883988298819880FFFFFFFFFFFFFFFF987F987E987D987C",
		x"98979896989598949893989298919890988F988E988D988C988B988A98899888",
		x"98A798A698A598A498A398A298A198A0989F989E989D989C989B989A98999898",
		x"98B798B698B598B498B398B298B198B098AF98AE98AD98AC98AB98AA98A998A8",
		x"98C398C298C198C0FFFFFFFFFFFFFFFF98BF98BE98BD98BC98BB98BA98B998B8",
		x"98D398D298D198D098CF98CE98CD98CC98CB98CA98C998C898C798C698C598C4",
		x"98E398E298E198E098DF98DE98DD98DC98DB98DA98D998D898D798D698D598D4",
		x"98F398F298F198F098EF98EE98ED98EC98EB98EA98E998E898E798E698E598E4",
		x"FFFFFFFFFFFFFFFF98FF98FE98FD98FC98FB98FA98F998F898F798F698F598F4",
		x"990F990E990D990C990B990A9909990899079906990599049903990299019900",
		x"991F991E991D991C991B991A9919991899179916991599149913991299119910",
		x"992F992E992D992C992B992A9929992899279926992599249923992299219920",
		x"993F993E993D993C993B993A9939993899379936993599349933993299319930",
		x"994B994A9949994899479946994599449943994299419940FFFFFFFFFFFFFFFF",
		x"995B995A9959995899579956995599549953995299519950994F994E994D994C",
		x"996B996A9969996899679966996599649963996299619960995F995E995D995C",
		x"997B997A9979997899779976997599749973997299719970996F996E996D996C",
		x"99879986998599849983998299819980FFFFFFFFFFFFFFFF997F997E997D997C",
		x"99979996999599949993999299919990998F998E998D998C998B998A99899988",
		x"99A799A699A599A499A399A299A199A0999F999E999D999C999B999A99999998",
		x"99B799B699B599B499B399B299B199B099AF99AE99AD99AC99AB99AA99A999A8",
		x"99C399C299C199C0FFFFFFFFFFFFFFFF99BF99BE99BD99BC99BB99BA99B999B8",
		x"99D399D299D199D099CF99CE99CD99CC99CB99CA99C999C899C799C699C599C4",
		x"99E399E299E199E099DF99DE99DD99DC99DB99DA99D999D899D799D699D599D4",
		x"99F399F299F199F099EF99EE99ED99EC99EB99EA99E999E899E799E699E599E4",
		x"FFFFFFFFFFFFFFFF99FF99FE99FD99FC99FB99FA99F999F899F799F699F599F4",
		x"9A0F9A0E9A0D9A0C9A0B9A0A9A099A089A079A069A059A049A039A029A019A00",
		x"9A1F9A1E9A1D9A1C9A1B9A1A9A199A189A179A169A159A149A139A129A119A10",
		x"9A2F9A2E9A2D9A2C9A2B9A2A9A299A289A279A269A259A249A239A229A219A20",
		x"9A3F9A3E9A3D9A3C9A3B9A3A9A399A389A379A369A359A349A339A329A319A30",
		x"9A4B9A4A9A499A489A479A469A459A449A439A429A419A40FFFFFFFFFFFFFFFF",
		x"9A5B9A5A9A599A589A579A569A559A549A539A529A519A509A4F9A4E9A4D9A4C",
		x"9A6B9A6A9A699A689A679A669A659A649A639A629A619A609A5F9A5E9A5D9A5C",
		x"9A7B9A7A9A799A789A779A769A759A749A739A729A719A709A6F9A6E9A6D9A6C",
		x"9A879A869A859A849A839A829A819A80FFFFFFFFFFFFFFFF9A7F9A7E9A7D9A7C",
		x"9A979A969A959A949A939A929A919A909A8F9A8E9A8D9A8C9A8B9A8A9A899A88",
		x"9AA79AA69AA59AA49AA39AA29AA19AA09A9F9A9E9A9D9A9C9A9B9A9A9A999A98",
		x"9AB79AB69AB59AB49AB39AB29AB19AB09AAF9AAE9AAD9AAC9AAB9AAA9AA99AA8",
		x"9AC39AC29AC19AC0FFFFFFFFFFFFFFFF9ABF9ABE9ABD9ABC9ABB9ABA9AB99AB8",
		x"9AD39AD29AD19AD09ACF9ACE9ACD9ACC9ACB9ACA9AC99AC89AC79AC69AC59AC4",
		x"9AE39AE29AE19AE09ADF9ADE9ADD9ADC9ADB9ADA9AD99AD89AD79AD69AD59AD4",
		x"9AF39AF29AF19AF09AEF9AEE9AED9AEC9AEB9AEA9AE99AE89AE79AE69AE59AE4",
		x"FFFFFFFFFFFFFFFF9AFF9AFE9AFD9AFC9AFB9AFA9AF99AF89AF79AF69AF59AF4",
		x"9B0F9B0E9B0D9B0C9B0B9B0A9B099B089B079B069B059B049B039B029B019B00",
		x"9B1F9B1E9B1D9B1C9B1B9B1A9B199B189B179B169B159B149B139B129B119B10",
		x"9B2F9B2E9B2D9B2C9B2B9B2A9B299B289B279B269B259B249B239B229B219B20",
		x"9B3F9B3E9B3D9B3C9B3B9B3A9B399B389B379B369B359B349B339B329B319B30",
		x"9B4B9B4A9B499B489B479B469B459B449B439B429B419B40FFFFFFFFFFFFFFFF",
		x"9B5B9B5A9B599B589B579B569B559B549B539B529B519B509B4F9B4E9B4D9B4C",
		x"9B6B9B6A9B699B689B679B669B659B649B639B629B619B609B5F9B5E9B5D9B5C",
		x"9B7B9B7A9B799B789B779B769B759B749B739B729B719B709B6F9B6E9B6D9B6C",
		x"9B879B869B859B849B839B829B819B80FFFFFFFFFFFFFFFF9B7F9B7E9B7D9B7C",
		x"9B979B969B959B949B939B929B919B909B8F9B8E9B8D9B8C9B8B9B8A9B899B88",
		x"9BA79BA69BA59BA49BA39BA29BA19BA09B9F9B9E9B9D9B9C9B9B9B9A9B999B98",
		x"9BB79BB69BB59BB49BB39BB29BB19BB09BAF9BAE9BAD9BAC9BAB9BAA9BA99BA8",
		x"9BC39BC29BC19BC0FFFFFFFFFFFFFFFF9BBF9BBE9BBD9BBC9BBB9BBA9BB99BB8",
		x"9BD39BD29BD19BD09BCF9BCE9BCD9BCC9BCB9BCA9BC99BC89BC79BC69BC59BC4",
		x"9BE39BE29BE19BE09BDF9BDE9BDD9BDC9BDB9BDA9BD99BD89BD79BD69BD59BD4",
		x"9BF39BF29BF19BF09BEF9BEE9BED9BEC9BEB9BEA9BE99BE89BE79BE69BE59BE4",
		x"FFFFFFFFFFFFFFFF9BFF9BFE9BFD9BFC9BFB9BFA9BF99BF89BF79BF69BF59BF4",
		x"9C0F9C0E9C0D9C0C9C0B9C0A9C099C089C079C069C059C049C039C029C019C00",
		x"9C1F9C1E9C1D9C1C9C1B9C1A9C199C189C179C169C159C149C139C129C119C10",
		x"9C2F9C2E9C2D9C2C9C2B9C2A9C299C289C279C269C259C249C239C229C219C20",
		x"9C3F9C3E9C3D9C3C9C3B9C3A9C399C389C379C369C359C349C339C329C319C30",
		x"9C4B9C4A9C499C489C479C469C459C449C439C429C419C40FFFFFFFFFFFFFFFF",
		x"9C5B9C5A9C599C589C579C569C559C549C539C529C519C509C4F9C4E9C4D9C4C",
		x"9C6B9C6A9C699C689C679C669C659C649C639C629C619C609C5F9C5E9C5D9C5C",
		x"9C7B9C7A9C799C789C779C769C759C749C739C729C719C709C6F9C6E9C6D9C6C",
		x"9C879C869C859C849C839C829C819C80FFFFFFFFFFFFFFFF9C7F9C7E9C7D9C7C",
		x"9C979C969C959C949C939C929C919C909C8F9C8E9C8D9C8C9C8B9C8A9C899C88",
		x"9CA79CA69CA59CA49CA39CA29CA19CA09C9F9C9E9C9D9C9C9C9B9C9A9C999C98",
		x"9CB79CB69CB59CB49CB39CB29CB19CB09CAF9CAE9CAD9CAC9CAB9CAA9CA99CA8",
		x"9CC39CC29CC19CC0FFFFFFFFFFFFFFFF9CBF9CBE9CBD9CBC9CBB9CBA9CB99CB8",
		x"9CD39CD29CD19CD09CCF9CCE9CCD9CCC9CCB9CCA9CC99CC89CC79CC69CC59CC4",
		x"9CE39CE29CE19CE09CDF9CDE9CDD9CDC9CDB9CDA9CD99CD89CD79CD69CD59CD4",
		x"9CF39CF29CF19CF09CEF9CEE9CED9CEC9CEB9CEA9CE99CE89CE79CE69CE59CE4",
		x"FFFFFFFFFFFFFFFF9CFF9CFE9CFD9CFC9CFB9CFA9CF99CF89CF79CF69CF59CF4",
		x"9D0F9D0E9D0D9D0C9D0B9D0A9D099D089D079D069D059D049D039D029D019D00",
		x"9D1F9D1E9D1D9D1C9D1B9D1A9D199D189D179D169D159D149D139D129D119D10",
		x"9D2F9D2E9D2D9D2C9D2B9D2A9D299D289D279D269D259D249D239D229D219D20",
		x"9D3F9D3E9D3D9D3C9D3B9D3A9D399D389D379D369D359D349D339D329D319D30",
		x"9D4B9D4A9D499D489D479D469D459D449D439D429D419D40FFFFFFFFFFFFFFFF",
		x"9D5B9D5A9D599D589D579D569D559D549D539D529D519D509D4F9D4E9D4D9D4C",
		x"9D6B9D6A9D699D689D679D669D659D649D639D629D619D609D5F9D5E9D5D9D5C",
		x"9D7B9D7A9D799D789D779D769D759D749D739D729D719D709D6F9D6E9D6D9D6C",
		x"9D879D869D859D849D839D829D819D80FFFFFFFFFFFFFFFF9D7F9D7E9D7D9D7C",
		x"9D979D969D959D949D939D929D919D909D8F9D8E9D8D9D8C9D8B9D8A9D899D88",
		x"9DA79DA69DA59DA49DA39DA29DA19DA09D9F9D9E9D9D9D9C9D9B9D9A9D999D98",
		x"9DB79DB69DB59DB49DB39DB29DB19DB09DAF9DAE9DAD9DAC9DAB9DAA9DA99DA8",
		x"9DC39DC29DC19DC0FFFFFFFFFFFFFFFF9DBF9DBE9DBD9DBC9DBB9DBA9DB99DB8",
		x"9DD39DD29DD19DD09DCF9DCE9DCD9DCC9DCB9DCA9DC99DC89DC79DC69DC59DC4",
		x"9DE39DE29DE19DE09DDF9DDE9DDD9DDC9DDB9DDA9DD99DD89DD79DD69DD59DD4",
		x"9DF39DF29DF19DF09DEF9DEE9DED9DEC9DEB9DEA9DE99DE89DE79DE69DE59DE4",
		x"FFFFFFFFFFFFFFFF9DFF9DFE9DFD9DFC9DFB9DFA9DF99DF89DF79DF69DF59DF4",
		x"9E0F9E0E9E0D9E0C9E0B9E0A9E099E089E079E069E059E049E039E029E019E00",
		x"9E1F9E1E9E1D9E1C9E1B9E1A9E199E189E179E169E159E149E139E129E119E10",
		x"9E2F9E2E9E2D9E2C9E2B9E2A9E299E289E279E269E259E249E239E229E219E20",
		x"9E3F9E3E9E3D9E3C9E3B9E3A9E399E389E379E369E359E349E339E329E319E30",
		x"9E4B9E4A9E499E489E479E469E459E449E439E429E419E40FFFFFFFFFFFFFFFF",
		x"9E5B9E5A9E599E589E579E569E559E549E539E529E519E509E4F9E4E9E4D9E4C",
		x"9E6B9E6A9E699E689E679E669E659E649E639E629E619E609E5F9E5E9E5D9E5C",
		x"9E7B9E7A9E799E789E779E769E759E749E739E729E719E709E6F9E6E9E6D9E6C",
		x"9E879E869E859E849E839E829E819E80FFFFFFFFFFFFFFFF9E7F9E7E9E7D9E7C",
		x"9E979E969E959E949E939E929E919E909E8F9E8E9E8D9E8C9E8B9E8A9E899E88",
		x"9EA79EA69EA59EA49EA39EA29EA19EA09E9F9E9E9E9D9E9C9E9B9E9A9E999E98",
		x"9EB79EB69EB59EB49EB39EB29EB19EB09EAF9EAE9EAD9EAC9EAB9EAA9EA99EA8",
		x"9EC39EC29EC19EC0FFFFFFFFFFFFFFFF9EBF9EBE9EBD9EBC9EBB9EBA9EB99EB8",
		x"9ED39ED29ED19ED09ECF9ECE9ECD9ECC9ECB9ECA9EC99EC89EC79EC69EC59EC4",
		x"9EE39EE29EE19EE09EDF9EDE9EDD9EDC9EDB9EDA9ED99ED89ED79ED69ED59ED4",
		x"9EF39EF29EF19EF09EEF9EEE9EED9EEC9EEB9EEA9EE99EE89EE79EE69EE59EE4",
		x"FFFFFFFFFFFFFFFF9EFF9EFE9EFD9EFC9EFB9EFA9EF99EF89EF79EF69EF59EF4",
		x"9F0F9F0E9F0D9F0C9F0B9F0A9F099F089F079F069F059F049F039F029F019F00",
		x"9F1F9F1E9F1D9F1C9F1B9F1A9F199F189F179F169F159F149F139F129F119F10",
		x"9F2F9F2E9F2D9F2C9F2B9F2A9F299F289F279F269F259F249F239F229F219F20",
		x"9F3F9F3E9F3D9F3C9F3B9F3A9F399F389F379F369F359F349F339F329F319F30",
		x"9F4B9F4A9F499F489F479F469F459F449F439F429F419F40FFFFFFFFFFFFFFFF",
		x"9F5B9F5A9F599F589F579F569F559F549F539F529F519F509F4F9F4E9F4D9F4C",
		x"9F6B9F6A9F699F689F679F669F659F649F639F629F619F609F5F9F5E9F5D9F5C",
		x"9F7B9F7A9F799F789F779F769F759F749F739F729F719F709F6F9F6E9F6D9F6C",
		x"9F879F869F859F849F839F829F819F80FFFFFFFFFFFFFFFF9F7F9F7E9F7D9F7C",
		x"9F979F969F959F949F939F929F919F909F8F9F8E9F8D9F8C9F8B9F8A9F899F88",
		x"9FA79FA69FA59FA49FA39FA29FA19FA09F9F9F9E9F9D9F9C9F9B9F9A9F999F98",
		x"9FB79FB69FB59FB49FB39FB29FB19FB09FAF9FAE9FAD9FAC9FAB9FAA9FA99FA8",
		x"9FC39FC29FC19FC0FFFFFFFFFFFFFFFF9FBF9FBE9FBD9FBC9FBB9FBA9FB99FB8",
		x"9FD39FD29FD19FD09FCF9FCE9FCD9FCC9FCB9FCA9FC99FC89FC79FC69FC59FC4",
		x"9FE39FE29FE19FE09FDF9FDE9FDD9FDC9FDB9FDA9FD99FD89FD79FD69FD59FD4",
		x"9FF39FF29FF19FF09FEF9FEE9FED9FEC9FEB9FEA9FE99FE89FE79FE69FE59FE4",
		x"FFFFFFFFFFFFFFFF9FFF9FFE9FFD9FFC9FFB9FFA9FF99FF89FF79FF69FF59FF4",
		x"A00FA00EA00DA00CA00BA00AA009A008A007A006A005A004A003A002A001A000",
		x"A01FA01EA01DA01CA01BA01AA019A018A017A016A015A014A013A012A011A010",
		x"A02FA02EA02DA02CA02BA02AA029A028A027A026A025A024A023A022A021A020",
		x"A03FA03EA03DA03CA03BA03AA039A038A037A036A035A034A033A032A031A030",
		x"A04BA04AA049A048A047A046A045A044A043A042A041A040FFFFFFFFFFFFFFFF",
		x"A05BA05AA059A058A057A056A055A054A053A052A051A050A04FA04EA04DA04C",
		x"A06BA06AA069A068A067A066A065A064A063A062A061A060A05FA05EA05DA05C",
		x"A07BA07AA079A078A077A076A075A074A073A072A071A070A06FA06EA06DA06C",
		x"A087A086A085A084A083A082A081A080FFFFFFFFFFFFFFFFA07FA07EA07DA07C",
		x"A097A096A095A094A093A092A091A090A08FA08EA08DA08CA08BA08AA089A088",
		x"A0A7A0A6A0A5A0A4A0A3A0A2A0A1A0A0A09FA09EA09DA09CA09BA09AA099A098",
		x"A0B7A0B6A0B5A0B4A0B3A0B2A0B1A0B0A0AFA0AEA0ADA0ACA0ABA0AAA0A9A0A8",
		x"A0C3A0C2A0C1A0C0FFFFFFFFFFFFFFFFA0BFA0BEA0BDA0BCA0BBA0BAA0B9A0B8",
		x"A0D3A0D2A0D1A0D0A0CFA0CEA0CDA0CCA0CBA0CAA0C9A0C8A0C7A0C6A0C5A0C4",
		x"A0E3A0E2A0E1A0E0A0DFA0DEA0DDA0DCA0DBA0DAA0D9A0D8A0D7A0D6A0D5A0D4",
		x"A0F3A0F2A0F1A0F0A0EFA0EEA0EDA0ECA0EBA0EAA0E9A0E8A0E7A0E6A0E5A0E4",
		x"FFFFFFFFFFFFFFFFA0FFA0FEA0FDA0FCA0FBA0FAA0F9A0F8A0F7A0F6A0F5A0F4",
		x"A10FA10EA10DA10CA10BA10AA109A108A107A106A105A104A103A102A101A100",
		x"A11FA11EA11DA11CA11BA11AA119A118A117A116A115A114A113A112A111A110",
		x"A12FA12EA12DA12CA12BA12AA129A128A127A126A125A124A123A122A121A120",
		x"A13FA13EA13DA13CA13BA13AA139A138A137A136A135A134A133A132A131A130",
		x"A14BA14AA149A148A147A146A145A144A143A142A141A140FFFFFFFFFFFFFFFF",
		x"A15BA15AA159A158A157A156A155A154A153A152A151A150A14FA14EA14DA14C",
		x"A16BA16AA169A168A167A166A165A164A163A162A161A160A15FA15EA15DA15C",
		x"A17BA17AA179A178A177A176A175A174A173A172A171A170A16FA16EA16DA16C",
		x"A187A186A185A184A183A182A181A180FFFFFFFFFFFFFFFFA17FA17EA17DA17C",
		x"A197A196A195A194A193A192A191A190A18FA18EA18DA18CA18BA18AA189A188",
		x"A1A7A1A6A1A5A1A4A1A3A1A2A1A1A1A0A19FA19EA19DA19CA19BA19AA199A198",
		x"A1B7A1B6A1B5A1B4A1B3A1B2A1B1A1B0A1AFA1AEA1ADA1ACA1ABA1AAA1A9A1A8",
		x"A1C3A1C2A1C1A1C0FFFFFFFFFFFFFFFFA1BFA1BEA1BDA1BCA1BBA1BAA1B9A1B8",
		x"A1D3A1D2A1D1A1D0A1CFA1CEA1CDA1CCA1CBA1CAA1C9A1C8A1C7A1C6A1C5A1C4",
		x"A1E3A1E2A1E1A1E0A1DFA1DEA1DDA1DCA1DBA1DAA1D9A1D8A1D7A1D6A1D5A1D4",
		x"A1F3A1F2A1F1A1F0A1EFA1EEA1EDA1ECA1EBA1EAA1E9A1E8A1E7A1E6A1E5A1E4",
		x"FFFFFFFFFFFFFFFFA1FFA1FEA1FDA1FCA1FBA1FAA1F9A1F8A1F7A1F6A1F5A1F4",
		x"A20FA20EA20DA20CA20BA20AA209A208A207A206A205A204A203A202A201A200",
		x"A21FA21EA21DA21CA21BA21AA219A218A217A216A215A214A213A212A211A210",
		x"A22FA22EA22DA22CA22BA22AA229A228A227A226A225A224A223A222A221A220",
		x"A23FA23EA23DA23CA23BA23AA239A238A237A236A235A234A233A232A231A230",
		x"A24BA24AA249A248A247A246A245A244A243A242A241A240FFFFFFFFFFFFFFFF",
		x"A25BA25AA259A258A257A256A255A254A253A252A251A250A24FA24EA24DA24C",
		x"A26BA26AA269A268A267A266A265A264A263A262A261A260A25FA25EA25DA25C",
		x"A27BA27AA279A278A277A276A275A274A273A272A271A270A26FA26EA26DA26C",
		x"A287A286A285A284A283A282A281A280FFFFFFFFFFFFFFFFA27FA27EA27DA27C",
		x"A297A296A295A294A293A292A291A290A28FA28EA28DA28CA28BA28AA289A288",
		x"A2A7A2A6A2A5A2A4A2A3A2A2A2A1A2A0A29FA29EA29DA29CA29BA29AA299A298",
		x"A2B7A2B6A2B5A2B4A2B3A2B2A2B1A2B0A2AFA2AEA2ADA2ACA2ABA2AAA2A9A2A8",
		x"A2C3A2C2A2C1A2C0FFFFFFFFFFFFFFFFA2BFA2BEA2BDA2BCA2BBA2BAA2B9A2B8",
		x"A2D3A2D2A2D1A2D0A2CFA2CEA2CDA2CCA2CBA2CAA2C9A2C8A2C7A2C6A2C5A2C4",
		x"A2E3A2E2A2E1A2E0A2DFA2DEA2DDA2DCA2DBA2DAA2D9A2D8A2D7A2D6A2D5A2D4",
		x"A2F3A2F2A2F1A2F0A2EFA2EEA2EDA2ECA2EBA2EAA2E9A2E8A2E7A2E6A2E5A2E4",
		x"FFFFFFFFFFFFFFFFA2FFA2FEA2FDA2FCA2FBA2FAA2F9A2F8A2F7A2F6A2F5A2F4",
		x"A30FA30EA30DA30CA30BA30AA309A308A307A306A305A304A303A302A301A300",
		x"A31FA31EA31DA31CA31BA31AA319A318A317A316A315A314A313A312A311A310",
		x"A32FA32EA32DA32CA32BA32AA329A328A327A326A325A324A323A322A321A320",
		x"A33FA33EA33DA33CA33BA33AA339A338A337A336A335A334A333A332A331A330",
		x"A34BA34AA349A348A347A346A345A344A343A342A341A340FFFFFFFFFFFFFFFF",
		x"A35BA35AA359A358A357A356A355A354A353A352A351A350A34FA34EA34DA34C",
		x"A36BA36AA369A368A367A366A365A364A363A362A361A360A35FA35EA35DA35C",
		x"A37BA37AA379A378A377A376A375A374A373A372A371A370A36FA36EA36DA36C",
		x"A387A386A385A384A383A382A381A380FFFFFFFFFFFFFFFFA37FA37EA37DA37C",
		x"A397A396A395A394A393A392A391A390A38FA38EA38DA38CA38BA38AA389A388",
		x"A3A7A3A6A3A5A3A4A3A3A3A2A3A1A3A0A39FA39EA39DA39CA39BA39AA399A398",
		x"A3B7A3B6A3B5A3B4A3B3A3B2A3B1A3B0A3AFA3AEA3ADA3ACA3ABA3AAA3A9A3A8",
		x"A3C3A3C2A3C1A3C0FFFFFFFFFFFFFFFFA3BFA3BEA3BDA3BCA3BBA3BAA3B9A3B8",
		x"A3D3A3D2A3D1A3D0A3CFA3CEA3CDA3CCA3CBA3CAA3C9A3C8A3C7A3C6A3C5A3C4",
		x"A3E3A3E2A3E1A3E0A3DFA3DEA3DDA3DCA3DBA3DAA3D9A3D8A3D7A3D6A3D5A3D4",
		x"A3F3A3F2A3F1A3F0A3EFA3EEA3EDA3ECA3EBA3EAA3E9A3E8A3E7A3E6A3E5A3E4",
		x"FFFFFFFFFFFFFFFFA3FFA3FEA3FDA3FCA3FBA3FAA3F9A3F8A3F7A3F6A3F5A3F4",
		x"A40FA40EA40DA40CA40BA40AA409A408A407A406A405A404A403A402A401A400",
		x"A41FA41EA41DA41CA41BA41AA419A418A417A416A415A414A413A412A411A410",
		x"A42FA42EA42DA42CA42BA42AA429A428A427A426A425A424A423A422A421A420",
		x"A43FA43EA43DA43CA43BA43AA439A438A437A436A435A434A433A432A431A430",
		x"A44BA44AA449A448A447A446A445A444A443A442A441A440FFFFFFFFFFFFFFFF",
		x"A45BA45AA459A458A457A456A455A454A453A452A451A450A44FA44EA44DA44C",
		x"A46BA46AA469A468A467A466A465A464A463A462A461A460A45FA45EA45DA45C",
		x"A47BA47AA479A478A477A476A475A474A473A472A471A470A46FA46EA46DA46C",
		x"A487A486A485A484A483A482A481A480FFFFFFFFFFFFFFFFA47FA47EA47DA47C",
		x"A497A496A495A494A493A492A491A490A48FA48EA48DA48CA48BA48AA489A488",
		x"A4A7A4A6A4A5A4A4A4A3A4A2A4A1A4A0A49FA49EA49DA49CA49BA49AA499A498",
		x"A4B7A4B6A4B5A4B4A4B3A4B2A4B1A4B0A4AFA4AEA4ADA4ACA4ABA4AAA4A9A4A8",
		x"A4C3A4C2A4C1A4C0FFFFFFFFFFFFFFFFA4BFA4BEA4BDA4BCA4BBA4BAA4B9A4B8",
		x"A4D3A4D2A4D1A4D0A4CFA4CEA4CDA4CCA4CBA4CAA4C9A4C8A4C7A4C6A4C5A4C4",
		x"A4E3A4E2A4E1A4E0A4DFA4DEA4DDA4DCA4DBA4DAA4D9A4D8A4D7A4D6A4D5A4D4",
		x"A4F3A4F2A4F1A4F0A4EFA4EEA4EDA4ECA4EBA4EAA4E9A4E8A4E7A4E6A4E5A4E4",
		x"FFFFFFFFFFFFFFFFA4FFA4FEA4FDA4FCA4FBA4FAA4F9A4F8A4F7A4F6A4F5A4F4",
		x"A50FA50EA50DA50CA50BA50AA509A508A507A506A505A504A503A502A501A500",
		x"A51FA51EA51DA51CA51BA51AA519A518A517A516A515A514A513A512A511A510",
		x"A52FA52EA52DA52CA52BA52AA529A528A527A526A525A524A523A522A521A520",
		x"A53FA53EA53DA53CA53BA53AA539A538A537A536A535A534A533A532A531A530",
		x"A54BA54AA549A548A547A546A545A544A543A542A541A540FFFFFFFFFFFFFFFF",
		x"A55BA55AA559A558A557A556A555A554A553A552A551A550A54FA54EA54DA54C",
		x"A56BA56AA569A568A567A566A565A564A563A562A561A560A55FA55EA55DA55C",
		x"A57BA57AA579A578A577A576A575A574A573A572A571A570A56FA56EA56DA56C",
		x"A587A586A585A584A583A582A581A580FFFFFFFFFFFFFFFFA57FA57EA57DA57C",
		x"A597A596A595A594A593A592A591A590A58FA58EA58DA58CA58BA58AA589A588",
		x"A5A7A5A6A5A5A5A4A5A3A5A2A5A1A5A0A59FA59EA59DA59CA59BA59AA599A598",
		x"A5B7A5B6A5B5A5B4A5B3A5B2A5B1A5B0A5AFA5AEA5ADA5ACA5ABA5AAA5A9A5A8",
		x"A5C3A5C2A5C1A5C0FFFFFFFFFFFFFFFFA5BFA5BEA5BDA5BCA5BBA5BAA5B9A5B8",
		x"A5D3A5D2A5D1A5D0A5CFA5CEA5CDA5CCA5CBA5CAA5C9A5C8A5C7A5C6A5C5A5C4",
		x"A5E3A5E2A5E1A5E0A5DFA5DEA5DDA5DCA5DBA5DAA5D9A5D8A5D7A5D6A5D5A5D4",
		x"A5F3A5F2A5F1A5F0A5EFA5EEA5EDA5ECA5EBA5EAA5E9A5E8A5E7A5E6A5E5A5E4",
		x"FFFFFFFFFFFFFFFFA5FFA5FEA5FDA5FCA5FBA5FAA5F9A5F8A5F7A5F6A5F5A5F4",
		x"A60FA60EA60DA60CA60BA60AA609A608A607A606A605A604A603A602A601A600",
		x"A61FA61EA61DA61CA61BA61AA619A618A617A616A615A614A613A612A611A610",
		x"A62FA62EA62DA62CA62BA62AA629A628A627A626A625A624A623A622A621A620",
		x"A63FA63EA63DA63CA63BA63AA639A638A637A636A635A634A633A632A631A630",
		x"A64BA64AA649A648A647A646A645A644A643A642A641A640FFFFFFFFFFFFFFFF",
		x"A65BA65AA659A658A657A656A655A654A653A652A651A650A64FA64EA64DA64C",
		x"A66BA66AA669A668A667A666A665A664A663A662A661A660A65FA65EA65DA65C",
		x"A67BA67AA679A678A677A676A675A674A673A672A671A670A66FA66EA66DA66C",
		x"A687A686A685A684A683A682A681A680FFFFFFFFFFFFFFFFA67FA67EA67DA67C",
		x"A697A696A695A694A693A692A691A690A68FA68EA68DA68CA68BA68AA689A688",
		x"A6A7A6A6A6A5A6A4A6A3A6A2A6A1A6A0A69FA69EA69DA69CA69BA69AA699A698",
		x"A6B7A6B6A6B5A6B4A6B3A6B2A6B1A6B0A6AFA6AEA6ADA6ACA6ABA6AAA6A9A6A8",
		x"A6C3A6C2A6C1A6C0FFFFFFFFFFFFFFFFA6BFA6BEA6BDA6BCA6BBA6BAA6B9A6B8",
		x"A6D3A6D2A6D1A6D0A6CFA6CEA6CDA6CCA6CBA6CAA6C9A6C8A6C7A6C6A6C5A6C4",
		x"A6E3A6E2A6E1A6E0A6DFA6DEA6DDA6DCA6DBA6DAA6D9A6D8A6D7A6D6A6D5A6D4",
		x"A6F3A6F2A6F1A6F0A6EFA6EEA6EDA6ECA6EBA6EAA6E9A6E8A6E7A6E6A6E5A6E4",
		x"FFFFFFFFFFFFFFFFA6FFA6FEA6FDA6FCA6FBA6FAA6F9A6F8A6F7A6F6A6F5A6F4",
		x"A70FA70EA70DA70CA70BA70AA709A708A707A706A705A704A703A702A701A700",
		x"A71FA71EA71DA71CA71BA71AA719A718A717A716A715A714A713A712A711A710",
		x"A72FA72EA72DA72CA72BA72AA729A728A727A726A725A724A723A722A721A720",
		x"A73FA73EA73DA73CA73BA73AA739A738A737A736A735A734A733A732A731A730",
		x"A74BA74AA749A748A747A746A745A744A743A742A741A740FFFFFFFFFFFFFFFF",
		x"A75BA75AA759A758A757A756A755A754A753A752A751A750A74FA74EA74DA74C",
		x"A76BA76AA769A768A767A766A765A764A763A762A761A760A75FA75EA75DA75C",
		x"A77BA77AA779A778A777A776A775A774A773A772A771A770A76FA76EA76DA76C",
		x"A787A786A785A784A783A782A781A780FFFFFFFFFFFFFFFFA77FA77EA77DA77C",
		x"A797A796A795A794A793A792A791A790A78FA78EA78DA78CA78BA78AA789A788",
		x"A7A7A7A6A7A5A7A4A7A3A7A2A7A1A7A0A79FA79EA79DA79CA79BA79AA799A798",
		x"A7B7A7B6A7B5A7B4A7B3A7B2A7B1A7B0A7AFA7AEA7ADA7ACA7ABA7AAA7A9A7A8",
		x"A7C3A7C2A7C1A7C0FFFFFFFFFFFFFFFFA7BFA7BEA7BDA7BCA7BBA7BAA7B9A7B8",
		x"A7D3A7D2A7D1A7D0A7CFA7CEA7CDA7CCA7CBA7CAA7C9A7C8A7C7A7C6A7C5A7C4",
		x"A7E3A7E2A7E1A7E0A7DFA7DEA7DDA7DCA7DBA7DAA7D9A7D8A7D7A7D6A7D5A7D4",
		x"A7F3A7F2A7F1A7F0A7EFA7EEA7EDA7ECA7EBA7EAA7E9A7E8A7E7A7E6A7E5A7E4",
		x"FFFFFFFFFFFFFFFFA7FFA7FEA7FDA7FCA7FBA7FAA7F9A7F8A7F7A7F6A7F5A7F4",
		x"A80FA80EA80DA80CA80BA80AA809A808A807A806A805A804A803A802A801A800",
		x"A81FA81EA81DA81CA81BA81AA819A818A817A816A815A814A813A812A811A810",
		x"A82FA82EA82DA82CA82BA82AA829A828A827A826A825A824A823A822A821A820",
		x"A83FA83EA83DA83CA83BA83AA839A838A837A836A835A834A833A832A831A830",
		x"A84BA84AA849A848A847A846A845A844A843A842A841A840FFFFFFFFFFFFFFFF",
		x"A85BA85AA859A858A857A856A855A854A853A852A851A850A84FA84EA84DA84C",
		x"A86BA86AA869A868A867A866A865A864A863A862A861A860A85FA85EA85DA85C",
		x"A87BA87AA879A878A877A876A875A874A873A872A871A870A86FA86EA86DA86C",
		x"A887A886A885A884A883A882A881A880FFFFFFFFFFFFFFFFA87FA87EA87DA87C",
		x"A897A896A895A894A893A892A891A890A88FA88EA88DA88CA88BA88AA889A888",
		x"A8A7A8A6A8A5A8A4A8A3A8A2A8A1A8A0A89FA89EA89DA89CA89BA89AA899A898",
		x"A8B7A8B6A8B5A8B4A8B3A8B2A8B1A8B0A8AFA8AEA8ADA8ACA8ABA8AAA8A9A8A8",
		x"A8C3A8C2A8C1A8C0FFFFFFFFFFFFFFFFA8BFA8BEA8BDA8BCA8BBA8BAA8B9A8B8",
		x"A8D3A8D2A8D1A8D0A8CFA8CEA8CDA8CCA8CBA8CAA8C9A8C8A8C7A8C6A8C5A8C4",
		x"A8E3A8E2A8E1A8E0A8DFA8DEA8DDA8DCA8DBA8DAA8D9A8D8A8D7A8D6A8D5A8D4",
		x"A8F3A8F2A8F1A8F0A8EFA8EEA8EDA8ECA8EBA8EAA8E9A8E8A8E7A8E6A8E5A8E4",
		x"FFFFFFFFFFFFFFFFA8FFA8FEA8FDA8FCA8FBA8FAA8F9A8F8A8F7A8F6A8F5A8F4",
		x"A90FA90EA90DA90CA90BA90AA909A908A907A906A905A904A903A902A901A900",
		x"A91FA91EA91DA91CA91BA91AA919A918A917A916A915A914A913A912A911A910",
		x"A92FA92EA92DA92CA92BA92AA929A928A927A926A925A924A923A922A921A920",
		x"A93FA93EA93DA93CA93BA93AA939A938A937A936A935A934A933A932A931A930",
		x"A94BA94AA949A948A947A946A945A944A943A942A941A940FFFFFFFFFFFFFFFF",
		x"A95BA95AA959A958A957A956A955A954A953A952A951A950A94FA94EA94DA94C",
		x"A96BA96AA969A968A967A966A965A964A963A962A961A960A95FA95EA95DA95C",
		x"A97BA97AA979A978A977A976A975A974A973A972A971A970A96FA96EA96DA96C",
		x"A987A986A985A984A983A982A981A980FFFFFFFFFFFFFFFFA97FA97EA97DA97C",
		x"A997A996A995A994A993A992A991A990A98FA98EA98DA98CA98BA98AA989A988",
		x"A9A7A9A6A9A5A9A4A9A3A9A2A9A1A9A0A99FA99EA99DA99CA99BA99AA999A998",
		x"A9B7A9B6A9B5A9B4A9B3A9B2A9B1A9B0A9AFA9AEA9ADA9ACA9ABA9AAA9A9A9A8",
		x"A9C3A9C2A9C1A9C0FFFFFFFFFFFFFFFFA9BFA9BEA9BDA9BCA9BBA9BAA9B9A9B8",
		x"A9D3A9D2A9D1A9D0A9CFA9CEA9CDA9CCA9CBA9CAA9C9A9C8A9C7A9C6A9C5A9C4",
		x"A9E3A9E2A9E1A9E0A9DFA9DEA9DDA9DCA9DBA9DAA9D9A9D8A9D7A9D6A9D5A9D4",
		x"A9F3A9F2A9F1A9F0A9EFA9EEA9EDA9ECA9EBA9EAA9E9A9E8A9E7A9E6A9E5A9E4",
		x"FFFFFFFFFFFFFFFFA9FFA9FEA9FDA9FCA9FBA9FAA9F9A9F8A9F7A9F6A9F5A9F4",
		x"AA0FAA0EAA0DAA0CAA0BAA0AAA09AA08AA07AA06AA05AA04AA03AA02AA01AA00",
		x"AA1FAA1EAA1DAA1CAA1BAA1AAA19AA18AA17AA16AA15AA14AA13AA12AA11AA10",
		x"AA2FAA2EAA2DAA2CAA2BAA2AAA29AA28AA27AA26AA25AA24AA23AA22AA21AA20",
		x"AA3FAA3EAA3DAA3CAA3BAA3AAA39AA38AA37AA36AA35AA34AA33AA32AA31AA30",
		x"AA4BAA4AAA49AA48AA47AA46AA45AA44AA43AA42AA41AA40FFFFFFFFFFFFFFFF",
		x"AA5BAA5AAA59AA58AA57AA56AA55AA54AA53AA52AA51AA50AA4FAA4EAA4DAA4C",
		x"AA6BAA6AAA69AA68AA67AA66AA65AA64AA63AA62AA61AA60AA5FAA5EAA5DAA5C",
		x"AA7BAA7AAA79AA78AA77AA76AA75AA74AA73AA72AA71AA70AA6FAA6EAA6DAA6C",
		x"AA87AA86AA85AA84AA83AA82AA81AA80FFFFFFFFFFFFFFFFAA7FAA7EAA7DAA7C",
		x"AA97AA96AA95AA94AA93AA92AA91AA90AA8FAA8EAA8DAA8CAA8BAA8AAA89AA88",
		x"AAA7AAA6AAA5AAA4AAA3AAA2AAA1AAA0AA9FAA9EAA9DAA9CAA9BAA9AAA99AA98",
		x"AAB7AAB6AAB5AAB4AAB3AAB2AAB1AAB0AAAFAAAEAAADAAACAAABAAAAAAA9AAA8",
		x"AAC3AAC2AAC1AAC0FFFFFFFFFFFFFFFFAABFAABEAABDAABCAABBAABAAAB9AAB8",
		x"AAD3AAD2AAD1AAD0AACFAACEAACDAACCAACBAACAAAC9AAC8AAC7AAC6AAC5AAC4",
		x"AAE3AAE2AAE1AAE0AADFAADEAADDAADCAADBAADAAAD9AAD8AAD7AAD6AAD5AAD4",
		x"AAF3AAF2AAF1AAF0AAEFAAEEAAEDAAECAAEBAAEAAAE9AAE8AAE7AAE6AAE5AAE4",
		x"FFFFFFFFFFFFFFFFAAFFAAFEAAFDAAFCAAFBAAFAAAF9AAF8AAF7AAF6AAF5AAF4",
		x"AB0FAB0EAB0DAB0CAB0BAB0AAB09AB08AB07AB06AB05AB04AB03AB02AB01AB00",
		x"AB1FAB1EAB1DAB1CAB1BAB1AAB19AB18AB17AB16AB15AB14AB13AB12AB11AB10",
		x"AB2FAB2EAB2DAB2CAB2BAB2AAB29AB28AB27AB26AB25AB24AB23AB22AB21AB20",
		x"AB3FAB3EAB3DAB3CAB3BAB3AAB39AB38AB37AB36AB35AB34AB33AB32AB31AB30",
		x"AB4BAB4AAB49AB48AB47AB46AB45AB44AB43AB42AB41AB40FFFFFFFFFFFFFFFF",
		x"AB5BAB5AAB59AB58AB57AB56AB55AB54AB53AB52AB51AB50AB4FAB4EAB4DAB4C",
		x"AB6BAB6AAB69AB68AB67AB66AB65AB64AB63AB62AB61AB60AB5FAB5EAB5DAB5C",
		x"AB7BAB7AAB79AB78AB77AB76AB75AB74AB73AB72AB71AB70AB6FAB6EAB6DAB6C",
		x"AB87AB86AB85AB84AB83AB82AB81AB80FFFFFFFFFFFFFFFFAB7FAB7EAB7DAB7C",
		x"AB97AB96AB95AB94AB93AB92AB91AB90AB8FAB8EAB8DAB8CAB8BAB8AAB89AB88",
		x"ABA7ABA6ABA5ABA4ABA3ABA2ABA1ABA0AB9FAB9EAB9DAB9CAB9BAB9AAB99AB98",
		x"ABB7ABB6ABB5ABB4ABB3ABB2ABB1ABB0ABAFABAEABADABACABABABAAABA9ABA8",
		x"ABC3ABC2ABC1ABC0FFFFFFFFFFFFFFFFABBFABBEABBDABBCABBBABBAABB9ABB8",
		x"ABD3ABD2ABD1ABD0ABCFABCEABCDABCCABCBABCAABC9ABC8ABC7ABC6ABC5ABC4",
		x"ABE3ABE2ABE1ABE0ABDFABDEABDDABDCABDBABDAABD9ABD8ABD7ABD6ABD5ABD4",
		x"ABF3ABF2ABF1ABF0ABEFABEEABEDABECABEBABEAABE9ABE8ABE7ABE6ABE5ABE4",
		x"FFFFFFFFFFFFFFFFABFFABFEABFDABFCABFBABFAABF9ABF8ABF7ABF6ABF5ABF4",
		x"AC0FAC0EAC0DAC0CAC0BAC0AAC09AC08AC07AC06AC05AC04AC03AC02AC01AC00",
		x"AC1FAC1EAC1DAC1CAC1BAC1AAC19AC18AC17AC16AC15AC14AC13AC12AC11AC10",
		x"AC2FAC2EAC2DAC2CAC2BAC2AAC29AC28AC27AC26AC25AC24AC23AC22AC21AC20",
		x"AC3FAC3EAC3DAC3CAC3BAC3AAC39AC38AC37AC36AC35AC34AC33AC32AC31AC30",
		x"AC4BAC4AAC49AC48AC47AC46AC45AC44AC43AC42AC41AC40FFFFFFFFFFFFFFFF",
		x"AC5BAC5AAC59AC58AC57AC56AC55AC54AC53AC52AC51AC50AC4FAC4EAC4DAC4C",
		x"AC6BAC6AAC69AC68AC67AC66AC65AC64AC63AC62AC61AC60AC5FAC5EAC5DAC5C",
		x"AC7BAC7AAC79AC78AC77AC76AC75AC74AC73AC72AC71AC70AC6FAC6EAC6DAC6C",
		x"AC87AC86AC85AC84AC83AC82AC81AC80FFFFFFFFFFFFFFFFAC7FAC7EAC7DAC7C",
		x"AC97AC96AC95AC94AC93AC92AC91AC90AC8FAC8EAC8DAC8CAC8BAC8AAC89AC88",
		x"ACA7ACA6ACA5ACA4ACA3ACA2ACA1ACA0AC9FAC9EAC9DAC9CAC9BAC9AAC99AC98",
		x"ACB7ACB6ACB5ACB4ACB3ACB2ACB1ACB0ACAFACAEACADACACACABACAAACA9ACA8",
		x"ACC3ACC2ACC1ACC0FFFFFFFFFFFFFFFFACBFACBEACBDACBCACBBACBAACB9ACB8",
		x"ACD3ACD2ACD1ACD0ACCFACCEACCDACCCACCBACCAACC9ACC8ACC7ACC6ACC5ACC4",
		x"ACE3ACE2ACE1ACE0ACDFACDEACDDACDCACDBACDAACD9ACD8ACD7ACD6ACD5ACD4",
		x"ACF3ACF2ACF1ACF0ACEFACEEACEDACECACEBACEAACE9ACE8ACE7ACE6ACE5ACE4",
		x"FFFFFFFFFFFFFFFFACFFACFEACFDACFCACFBACFAACF9ACF8ACF7ACF6ACF5ACF4",
		x"AD0FAD0EAD0DAD0CAD0BAD0AAD09AD08AD07AD06AD05AD04AD03AD02AD01AD00",
		x"AD1FAD1EAD1DAD1CAD1BAD1AAD19AD18AD17AD16AD15AD14AD13AD12AD11AD10",
		x"AD2FAD2EAD2DAD2CAD2BAD2AAD29AD28AD27AD26AD25AD24AD23AD22AD21AD20",
		x"AD3FAD3EAD3DAD3CAD3BAD3AAD39AD38AD37AD36AD35AD34AD33AD32AD31AD30",
		x"AD4BAD4AAD49AD48AD47AD46AD45AD44AD43AD42AD41AD40FFFFFFFFFFFFFFFF",
		x"AD5BAD5AAD59AD58AD57AD56AD55AD54AD53AD52AD51AD50AD4FAD4EAD4DAD4C",
		x"AD6BAD6AAD69AD68AD67AD66AD65AD64AD63AD62AD61AD60AD5FAD5EAD5DAD5C",
		x"AD7BAD7AAD79AD78AD77AD76AD75AD74AD73AD72AD71AD70AD6FAD6EAD6DAD6C",
		x"AD87AD86AD85AD84AD83AD82AD81AD80FFFFFFFFFFFFFFFFAD7FAD7EAD7DAD7C",
		x"AD97AD96AD95AD94AD93AD92AD91AD90AD8FAD8EAD8DAD8CAD8BAD8AAD89AD88",
		x"ADA7ADA6ADA5ADA4ADA3ADA2ADA1ADA0AD9FAD9EAD9DAD9CAD9BAD9AAD99AD98",
		x"ADB7ADB6ADB5ADB4ADB3ADB2ADB1ADB0ADAFADAEADADADACADABADAAADA9ADA8",
		x"ADC3ADC2ADC1ADC0FFFFFFFFFFFFFFFFADBFADBEADBDADBCADBBADBAADB9ADB8",
		x"ADD3ADD2ADD1ADD0ADCFADCEADCDADCCADCBADCAADC9ADC8ADC7ADC6ADC5ADC4",
		x"ADE3ADE2ADE1ADE0ADDFADDEADDDADDCADDBADDAADD9ADD8ADD7ADD6ADD5ADD4",
		x"ADF3ADF2ADF1ADF0ADEFADEEADEDADECADEBADEAADE9ADE8ADE7ADE6ADE5ADE4",
		x"FFFFFFFFFFFFFFFFADFFADFEADFDADFCADFBADFAADF9ADF8ADF7ADF6ADF5ADF4",
		x"AE0FAE0EAE0DAE0CAE0BAE0AAE09AE08AE07AE06AE05AE04AE03AE02AE01AE00",
		x"AE1FAE1EAE1DAE1CAE1BAE1AAE19AE18AE17AE16AE15AE14AE13AE12AE11AE10",
		x"AE2FAE2EAE2DAE2CAE2BAE2AAE29AE28AE27AE26AE25AE24AE23AE22AE21AE20",
		x"AE3FAE3EAE3DAE3CAE3BAE3AAE39AE38AE37AE36AE35AE34AE33AE32AE31AE30",
		x"AE4BAE4AAE49AE48AE47AE46AE45AE44AE43AE42AE41AE40FFFFFFFFFFFFFFFF",
		x"AE5BAE5AAE59AE58AE57AE56AE55AE54AE53AE52AE51AE50AE4FAE4EAE4DAE4C",
		x"AE6BAE6AAE69AE68AE67AE66AE65AE64AE63AE62AE61AE60AE5FAE5EAE5DAE5C",
		x"AE7BAE7AAE79AE78AE77AE76AE75AE74AE73AE72AE71AE70AE6FAE6EAE6DAE6C",
		x"AE87AE86AE85AE84AE83AE82AE81AE80FFFFFFFFFFFFFFFFAE7FAE7EAE7DAE7C",
		x"AE97AE96AE95AE94AE93AE92AE91AE90AE8FAE8EAE8DAE8CAE8BAE8AAE89AE88",
		x"AEA7AEA6AEA5AEA4AEA3AEA2AEA1AEA0AE9FAE9EAE9DAE9CAE9BAE9AAE99AE98",
		x"AEB7AEB6AEB5AEB4AEB3AEB2AEB1AEB0AEAFAEAEAEADAEACAEABAEAAAEA9AEA8",
		x"AEC3AEC2AEC1AEC0FFFFFFFFFFFFFFFFAEBFAEBEAEBDAEBCAEBBAEBAAEB9AEB8",
		x"AED3AED2AED1AED0AECFAECEAECDAECCAECBAECAAEC9AEC8AEC7AEC6AEC5AEC4",
		x"AEE3AEE2AEE1AEE0AEDFAEDEAEDDAEDCAEDBAEDAAED9AED8AED7AED6AED5AED4",
		x"AEF3AEF2AEF1AEF0AEEFAEEEAEEDAEECAEEBAEEAAEE9AEE8AEE7AEE6AEE5AEE4",
		x"FFFFFFFFFFFFFFFFAEFFAEFEAEFDAEFCAEFBAEFAAEF9AEF8AEF7AEF6AEF5AEF4",
		x"AF0FAF0EAF0DAF0CAF0BAF0AAF09AF08AF07AF06AF05AF04AF03AF02AF01AF00",
		x"AF1FAF1EAF1DAF1CAF1BAF1AAF19AF18AF17AF16AF15AF14AF13AF12AF11AF10",
		x"AF2FAF2EAF2DAF2CAF2BAF2AAF29AF28AF27AF26AF25AF24AF23AF22AF21AF20",
		x"AF3FAF3EAF3DAF3CAF3BAF3AAF39AF38AF37AF36AF35AF34AF33AF32AF31AF30",
		x"AF4BAF4AAF49AF48AF47AF46AF45AF44AF43AF42AF41AF40FFFFFFFFFFFFFFFF",
		x"AF5BAF5AAF59AF58AF57AF56AF55AF54AF53AF52AF51AF50AF4FAF4EAF4DAF4C",
		x"AF6BAF6AAF69AF68AF67AF66AF65AF64AF63AF62AF61AF60AF5FAF5EAF5DAF5C",
		x"AF7BAF7AAF79AF78AF77AF76AF75AF74AF73AF72AF71AF70AF6FAF6EAF6DAF6C",
		x"AF87AF86AF85AF84AF83AF82AF81AF80FFFFFFFFFFFFFFFFAF7FAF7EAF7DAF7C",
		x"AF97AF96AF95AF94AF93AF92AF91AF90AF8FAF8EAF8DAF8CAF8BAF8AAF89AF88",
		x"AFA7AFA6AFA5AFA4AFA3AFA2AFA1AFA0AF9FAF9EAF9DAF9CAF9BAF9AAF99AF98",
		x"AFB7AFB6AFB5AFB4AFB3AFB2AFB1AFB0AFAFAFAEAFADAFACAFABAFAAAFA9AFA8",
		x"AFC3AFC2AFC1AFC0FFFFFFFFFFFFFFFFAFBFAFBEAFBDAFBCAFBBAFBAAFB9AFB8",
		x"AFD3AFD2AFD1AFD0AFCFAFCEAFCDAFCCAFCBAFCAAFC9AFC8AFC7AFC6AFC5AFC4",
		x"AFE3AFE2AFE1AFE0AFDFAFDEAFDDAFDCAFDBAFDAAFD9AFD8AFD7AFD6AFD5AFD4",
		x"AFF3AFF2AFF1AFF0AFEFAFEEAFEDAFECAFEBAFEAAFE9AFE8AFE7AFE6AFE5AFE4",
		x"FFFFFFFFFFFFFFFFAFFFAFFEAFFDAFFCAFFBAFFAAFF9AFF8AFF7AFF6AFF5AFF4",
		x"B00FB00EB00DB00CB00BB00AB009B008B007B006B005B004B003B002B001B000",
		x"B01FB01EB01DB01CB01BB01AB019B018B017B016B015B014B013B012B011B010",
		x"B02FB02EB02DB02CB02BB02AB029B028B027B026B025B024B023B022B021B020",
		x"B03FB03EB03DB03CB03BB03AB039B038B037B036B035B034B033B032B031B030",
		x"B04BB04AB049B048B047B046B045B044B043B042B041B040FFFFFFFFFFFFFFFF",
		x"B05BB05AB059B058B057B056B055B054B053B052B051B050B04FB04EB04DB04C",
		x"B06BB06AB069B068B067B066B065B064B063B062B061B060B05FB05EB05DB05C",
		x"B07BB07AB079B078B077B076B075B074B073B072B071B070B06FB06EB06DB06C",
		x"B087B086B085B084B083B082B081B080FFFFFFFFFFFFFFFFB07FB07EB07DB07C",
		x"B097B096B095B094B093B092B091B090B08FB08EB08DB08CB08BB08AB089B088",
		x"B0A7B0A6B0A5B0A4B0A3B0A2B0A1B0A0B09FB09EB09DB09CB09BB09AB099B098",
		x"B0B7B0B6B0B5B0B4B0B3B0B2B0B1B0B0B0AFB0AEB0ADB0ACB0ABB0AAB0A9B0A8",
		x"B0C3B0C2B0C1B0C0FFFFFFFFFFFFFFFFB0BFB0BEB0BDB0BCB0BBB0BAB0B9B0B8",
		x"B0D3B0D2B0D1B0D0B0CFB0CEB0CDB0CCB0CBB0CAB0C9B0C8B0C7B0C6B0C5B0C4",
		x"B0E3B0E2B0E1B0E0B0DFB0DEB0DDB0DCB0DBB0DAB0D9B0D8B0D7B0D6B0D5B0D4",
		x"B0F3B0F2B0F1B0F0B0EFB0EEB0EDB0ECB0EBB0EAB0E9B0E8B0E7B0E6B0E5B0E4",
		x"FFFFFFFFFFFFFFFFB0FFB0FEB0FDB0FCB0FBB0FAB0F9B0F8B0F7B0F6B0F5B0F4",
		x"B10FB10EB10DB10CB10BB10AB109B108B107B106B105B104B103B102B101B100",
		x"B11FB11EB11DB11CB11BB11AB119B118B117B116B115B114B113B112B111B110",
		x"B12FB12EB12DB12CB12BB12AB129B128B127B126B125B124B123B122B121B120",
		x"B13FB13EB13DB13CB13BB13AB139B138B137B136B135B134B133B132B131B130",
		x"B14BB14AB149B148B147B146B145B144B143B142B141B140FFFFFFFFFFFFFFFF",
		x"B15BB15AB159B158B157B156B155B154B153B152B151B150B14FB14EB14DB14C",
		x"B16BB16AB169B168B167B166B165B164B163B162B161B160B15FB15EB15DB15C",
		x"B17BB17AB179B178B177B176B175B174B173B172B171B170B16FB16EB16DB16C",
		x"B187B186B185B184B183B182B181B180FFFFFFFFFFFFFFFFB17FB17EB17DB17C",
		x"B197B196B195B194B193B192B191B190B18FB18EB18DB18CB18BB18AB189B188",
		x"B1A7B1A6B1A5B1A4B1A3B1A2B1A1B1A0B19FB19EB19DB19CB19BB19AB199B198",
		x"B1B7B1B6B1B5B1B4B1B3B1B2B1B1B1B0B1AFB1AEB1ADB1ACB1ABB1AAB1A9B1A8",
		x"B1C3B1C2B1C1B1C0FFFFFFFFFFFFFFFFB1BFB1BEB1BDB1BCB1BBB1BAB1B9B1B8",
		x"B1D3B1D2B1D1B1D0B1CFB1CEB1CDB1CCB1CBB1CAB1C9B1C8B1C7B1C6B1C5B1C4",
		x"B1E3B1E2B1E1B1E0B1DFB1DEB1DDB1DCB1DBB1DAB1D9B1D8B1D7B1D6B1D5B1D4",
		x"B1F3B1F2B1F1B1F0B1EFB1EEB1EDB1ECB1EBB1EAB1E9B1E8B1E7B1E6B1E5B1E4",
		x"FFFFFFFFFFFFFFFFB1FFB1FEB1FDB1FCB1FBB1FAB1F9B1F8B1F7B1F6B1F5B1F4",
		x"B20FB20EB20DB20CB20BB20AB209B208B207B206B205B204B203B202B201B200",
		x"B21FB21EB21DB21CB21BB21AB219B218B217B216B215B214B213B212B211B210",
		x"B22FB22EB22DB22CB22BB22AB229B228B227B226B225B224B223B222B221B220",
		x"B23FB23EB23DB23CB23BB23AB239B238B237B236B235B234B233B232B231B230",
		x"B24BB24AB249B248B247B246B245B244B243B242B241B240FFFFFFFFFFFFFFFF",
		x"B25BB25AB259B258B257B256B255B254B253B252B251B250B24FB24EB24DB24C",
		x"B26BB26AB269B268B267B266B265B264B263B262B261B260B25FB25EB25DB25C",
		x"B27BB27AB279B278B277B276B275B274B273B272B271B270B26FB26EB26DB26C",
		x"B287B286B285B284B283B282B281B280FFFFFFFFFFFFFFFFB27FB27EB27DB27C",
		x"B297B296B295B294B293B292B291B290B28FB28EB28DB28CB28BB28AB289B288",
		x"B2A7B2A6B2A5B2A4B2A3B2A2B2A1B2A0B29FB29EB29DB29CB29BB29AB299B298",
		x"B2B7B2B6B2B5B2B4B2B3B2B2B2B1B2B0B2AFB2AEB2ADB2ACB2ABB2AAB2A9B2A8",
		x"B2C3B2C2B2C1B2C0FFFFFFFFFFFFFFFFB2BFB2BEB2BDB2BCB2BBB2BAB2B9B2B8",
		x"B2D3B2D2B2D1B2D0B2CFB2CEB2CDB2CCB2CBB2CAB2C9B2C8B2C7B2C6B2C5B2C4",
		x"B2E3B2E2B2E1B2E0B2DFB2DEB2DDB2DCB2DBB2DAB2D9B2D8B2D7B2D6B2D5B2D4",
		x"B2F3B2F2B2F1B2F0B2EFB2EEB2EDB2ECB2EBB2EAB2E9B2E8B2E7B2E6B2E5B2E4",
		x"FFFFFFFFFFFFFFFFB2FFB2FEB2FDB2FCB2FBB2FAB2F9B2F8B2F7B2F6B2F5B2F4",
		x"B30FB30EB30DB30CB30BB30AB309B308B307B306B305B304B303B302B301B300",
		x"B31FB31EB31DB31CB31BB31AB319B318B317B316B315B314B313B312B311B310",
		x"B32FB32EB32DB32CB32BB32AB329B328B327B326B325B324B323B322B321B320",
		x"B33FB33EB33DB33CB33BB33AB339B338B337B336B335B334B333B332B331B330",
		x"B34BB34AB349B348B347B346B345B344B343B342B341B340FFFFFFFFFFFFFFFF",
		x"B35BB35AB359B358B357B356B355B354B353B352B351B350B34FB34EB34DB34C",
		x"B36BB36AB369B368B367B366B365B364B363B362B361B360B35FB35EB35DB35C",
		x"B37BB37AB379B378B377B376B375B374B373B372B371B370B36FB36EB36DB36C",
		x"B387B386B385B384B383B382B381B380FFFFFFFFFFFFFFFFB37FB37EB37DB37C",
		x"B397B396B395B394B393B392B391B390B38FB38EB38DB38CB38BB38AB389B388",
		x"B3A7B3A6B3A5B3A4B3A3B3A2B3A1B3A0B39FB39EB39DB39CB39BB39AB399B398",
		x"B3B7B3B6B3B5B3B4B3B3B3B2B3B1B3B0B3AFB3AEB3ADB3ACB3ABB3AAB3A9B3A8",
		x"B3C3B3C2B3C1B3C0FFFFFFFFFFFFFFFFB3BFB3BEB3BDB3BCB3BBB3BAB3B9B3B8",
		x"B3D3B3D2B3D1B3D0B3CFB3CEB3CDB3CCB3CBB3CAB3C9B3C8B3C7B3C6B3C5B3C4",
		x"B3E3B3E2B3E1B3E0B3DFB3DEB3DDB3DCB3DBB3DAB3D9B3D8B3D7B3D6B3D5B3D4",
		x"B3F3B3F2B3F1B3F0B3EFB3EEB3EDB3ECB3EBB3EAB3E9B3E8B3E7B3E6B3E5B3E4",
		x"FFFFFFFFFFFFFFFFB3FFB3FEB3FDB3FCB3FBB3FAB3F9B3F8B3F7B3F6B3F5B3F4",
		x"B40FB40EB40DB40CB40BB40AB409B408B407B406B405B404B403B402B401B400",
		x"B41FB41EB41DB41CB41BB41AB419B418B417B416B415B414B413B412B411B410",
		x"B42FB42EB42DB42CB42BB42AB429B428B427B426B425B424B423B422B421B420",
		x"B43FB43EB43DB43CB43BB43AB439B438B437B436B435B434B433B432B431B430",
		x"B44BB44AB449B448B447B446B445B444B443B442B441B440FFFFFFFFFFFFFFFF",
		x"B45BB45AB459B458B457B456B455B454B453B452B451B450B44FB44EB44DB44C",
		x"B46BB46AB469B468B467B466B465B464B463B462B461B460B45FB45EB45DB45C",
		x"B47BB47AB479B478B477B476B475B474B473B472B471B470B46FB46EB46DB46C",
		x"B487B486B485B484B483B482B481B480FFFFFFFFFFFFFFFFB47FB47EB47DB47C",
		x"B497B496B495B494B493B492B491B490B48FB48EB48DB48CB48BB48AB489B488",
		x"B4A7B4A6B4A5B4A4B4A3B4A2B4A1B4A0B49FB49EB49DB49CB49BB49AB499B498",
		x"B4B7B4B6B4B5B4B4B4B3B4B2B4B1B4B0B4AFB4AEB4ADB4ACB4ABB4AAB4A9B4A8",
		x"B4C3B4C2B4C1B4C0FFFFFFFFFFFFFFFFB4BFB4BEB4BDB4BCB4BBB4BAB4B9B4B8",
		x"B4D3B4D2B4D1B4D0B4CFB4CEB4CDB4CCB4CBB4CAB4C9B4C8B4C7B4C6B4C5B4C4",
		x"B4E3B4E2B4E1B4E0B4DFB4DEB4DDB4DCB4DBB4DAB4D9B4D8B4D7B4D6B4D5B4D4",
		x"B4F3B4F2B4F1B4F0B4EFB4EEB4EDB4ECB4EBB4EAB4E9B4E8B4E7B4E6B4E5B4E4",
		x"FFFFFFFFFFFFFFFFB4FFB4FEB4FDB4FCB4FBB4FAB4F9B4F8B4F7B4F6B4F5B4F4",
		x"B50FB50EB50DB50CB50BB50AB509B508B507B506B505B504B503B502B501B500",
		x"B51FB51EB51DB51CB51BB51AB519B518B517B516B515B514B513B512B511B510",
		x"B52FB52EB52DB52CB52BB52AB529B528B527B526B525B524B523B522B521B520",
		x"B53FB53EB53DB53CB53BB53AB539B538B537B536B535B534B533B532B531B530",
		x"B54BB54AB549B548B547B546B545B544B543B542B541B540FFFFFFFFFFFFFFFF",
		x"B55BB55AB559B558B557B556B555B554B553B552B551B550B54FB54EB54DB54C",
		x"B56BB56AB569B568B567B566B565B564B563B562B561B560B55FB55EB55DB55C",
		x"B57BB57AB579B578B577B576B575B574B573B572B571B570B56FB56EB56DB56C",
		x"B587B586B585B584B583B582B581B580FFFFFFFFFFFFFFFFB57FB57EB57DB57C",
		x"B597B596B595B594B593B592B591B590B58FB58EB58DB58CB58BB58AB589B588",
		x"B5A7B5A6B5A5B5A4B5A3B5A2B5A1B5A0B59FB59EB59DB59CB59BB59AB599B598",
		x"B5B7B5B6B5B5B5B4B5B3B5B2B5B1B5B0B5AFB5AEB5ADB5ACB5ABB5AAB5A9B5A8",
		x"B5C3B5C2B5C1B5C0FFFFFFFFFFFFFFFFB5BFB5BEB5BDB5BCB5BBB5BAB5B9B5B8",
		x"B5D3B5D2B5D1B5D0B5CFB5CEB5CDB5CCB5CBB5CAB5C9B5C8B5C7B5C6B5C5B5C4",
		x"B5E3B5E2B5E1B5E0B5DFB5DEB5DDB5DCB5DBB5DAB5D9B5D8B5D7B5D6B5D5B5D4",
		x"B5F3B5F2B5F1B5F0B5EFB5EEB5EDB5ECB5EBB5EAB5E9B5E8B5E7B5E6B5E5B5E4",
		x"FFFFFFFFFFFFFFFFB5FFB5FEB5FDB5FCB5FBB5FAB5F9B5F8B5F7B5F6B5F5B5F4",
		x"B60FB60EB60DB60CB60BB60AB609B608B607B606B605B604B603B602B601B600",
		x"B61FB61EB61DB61CB61BB61AB619B618B617B616B615B614B613B612B611B610",
		x"B62FB62EB62DB62CB62BB62AB629B628B627B626B625B624B623B622B621B620",
		x"B63FB63EB63DB63CB63BB63AB639B638B637B636B635B634B633B632B631B630",
		x"B64BB64AB649B648B647B646B645B644B643B642B641B640FFFFFFFFFFFFFFFF",
		x"B65BB65AB659B658B657B656B655B654B653B652B651B650B64FB64EB64DB64C",
		x"B66BB66AB669B668B667B666B665B664B663B662B661B660B65FB65EB65DB65C",
		x"B67BB67AB679B678B677B676B675B674B673B672B671B670B66FB66EB66DB66C",
		x"B687B686B685B684B683B682B681B680FFFFFFFFFFFFFFFFB67FB67EB67DB67C",
		x"B697B696B695B694B693B692B691B690B68FB68EB68DB68CB68BB68AB689B688",
		x"B6A7B6A6B6A5B6A4B6A3B6A2B6A1B6A0B69FB69EB69DB69CB69BB69AB699B698",
		x"B6B7B6B6B6B5B6B4B6B3B6B2B6B1B6B0B6AFB6AEB6ADB6ACB6ABB6AAB6A9B6A8",
		x"B6C3B6C2B6C1B6C0FFFFFFFFFFFFFFFFB6BFB6BEB6BDB6BCB6BBB6BAB6B9B6B8",
		x"B6D3B6D2B6D1B6D0B6CFB6CEB6CDB6CCB6CBB6CAB6C9B6C8B6C7B6C6B6C5B6C4",
		x"B6E3B6E2B6E1B6E0B6DFB6DEB6DDB6DCB6DBB6DAB6D9B6D8B6D7B6D6B6D5B6D4",
		x"B6F3B6F2B6F1B6F0B6EFB6EEB6EDB6ECB6EBB6EAB6E9B6E8B6E7B6E6B6E5B6E4",
		x"FFFFFFFFFFFFFFFFB6FFB6FEB6FDB6FCB6FBB6FAB6F9B6F8B6F7B6F6B6F5B6F4",
		x"B70FB70EB70DB70CB70BB70AB709B708B707B706B705B704B703B702B701B700",
		x"B71FB71EB71DB71CB71BB71AB719B718B717B716B715B714B713B712B711B710",
		x"B72FB72EB72DB72CB72BB72AB729B728B727B726B725B724B723B722B721B720",
		x"B73FB73EB73DB73CB73BB73AB739B738B737B736B735B734B733B732B731B730",
		x"B74BB74AB749B748B747B746B745B744B743B742B741B740FFFFFFFFFFFFFFFF",
		x"B75BB75AB759B758B757B756B755B754B753B752B751B750B74FB74EB74DB74C",
		x"B76BB76AB769B768B767B766B765B764B763B762B761B760B75FB75EB75DB75C",
		x"B77BB77AB779B778B777B776B775B774B773B772B771B770B76FB76EB76DB76C",
		x"B787B786B785B784B783B782B781B780FFFFFFFFFFFFFFFFB77FB77EB77DB77C",
		x"B797B796B795B794B793B792B791B790B78FB78EB78DB78CB78BB78AB789B788",
		x"B7A7B7A6B7A5B7A4B7A3B7A2B7A1B7A0B79FB79EB79DB79CB79BB79AB799B798",
		x"B7B7B7B6B7B5B7B4B7B3B7B2B7B1B7B0B7AFB7AEB7ADB7ACB7ABB7AAB7A9B7A8",
		x"B7C3B7C2B7C1B7C0FFFFFFFFFFFFFFFFB7BFB7BEB7BDB7BCB7BBB7BAB7B9B7B8",
		x"B7D3B7D2B7D1B7D0B7CFB7CEB7CDB7CCB7CBB7CAB7C9B7C8B7C7B7C6B7C5B7C4",
		x"B7E3B7E2B7E1B7E0B7DFB7DEB7DDB7DCB7DBB7DAB7D9B7D8B7D7B7D6B7D5B7D4",
		x"B7F3B7F2B7F1B7F0B7EFB7EEB7EDB7ECB7EBB7EAB7E9B7E8B7E7B7E6B7E5B7E4",
		x"FFFFFFFFFFFFFFFFB7FFB7FEB7FDB7FCB7FBB7FAB7F9B7F8B7F7B7F6B7F5B7F4",
		x"B80FB80EB80DB80CB80BB80AB809B808B807B806B805B804B803B802B801B800",
		x"B81FB81EB81DB81CB81BB81AB819B818B817B816B815B814B813B812B811B810",
		x"B82FB82EB82DB82CB82BB82AB829B828B827B826B825B824B823B822B821B820",
		x"B83FB83EB83DB83CB83BB83AB839B838B837B836B835B834B833B832B831B830",
		x"B84BB84AB849B848B847B846B845B844B843B842B841B840FFFFFFFFFFFFFFFF",
		x"B85BB85AB859B858B857B856B855B854B853B852B851B850B84FB84EB84DB84C",
		x"B86BB86AB869B868B867B866B865B864B863B862B861B860B85FB85EB85DB85C",
		x"B87BB87AB879B878B877B876B875B874B873B872B871B870B86FB86EB86DB86C",
		x"B887B886B885B884B883B882B881B880FFFFFFFFFFFFFFFFB87FB87EB87DB87C",
		x"B897B896B895B894B893B892B891B890B88FB88EB88DB88CB88BB88AB889B888",
		x"B8A7B8A6B8A5B8A4B8A3B8A2B8A1B8A0B89FB89EB89DB89CB89BB89AB899B898",
		x"B8B7B8B6B8B5B8B4B8B3B8B2B8B1B8B0B8AFB8AEB8ADB8ACB8ABB8AAB8A9B8A8",
		x"B8C3B8C2B8C1B8C0FFFFFFFFFFFFFFFFB8BFB8BEB8BDB8BCB8BBB8BAB8B9B8B8",
		x"B8D3B8D2B8D1B8D0B8CFB8CEB8CDB8CCB8CBB8CAB8C9B8C8B8C7B8C6B8C5B8C4",
		x"B8E3B8E2B8E1B8E0B8DFB8DEB8DDB8DCB8DBB8DAB8D9B8D8B8D7B8D6B8D5B8D4",
		x"B8F3B8F2B8F1B8F0B8EFB8EEB8EDB8ECB8EBB8EAB8E9B8E8B8E7B8E6B8E5B8E4",
		x"FFFFFFFFFFFFFFFFB8FFB8FEB8FDB8FCB8FBB8FAB8F9B8F8B8F7B8F6B8F5B8F4",
		x"B90FB90EB90DB90CB90BB90AB909B908B907B906B905B904B903B902B901B900",
		x"B91FB91EB91DB91CB91BB91AB919B918B917B916B915B914B913B912B911B910",
		x"B92FB92EB92DB92CB92BB92AB929B928B927B926B925B924B923B922B921B920",
		x"B93FB93EB93DB93CB93BB93AB939B938B937B936B935B934B933B932B931B930",
		x"B94BB94AB949B948B947B946B945B944B943B942B941B940FFFFFFFFFFFFFFFF",
		x"B95BB95AB959B958B957B956B955B954B953B952B951B950B94FB94EB94DB94C",
		x"B96BB96AB969B968B967B966B965B964B963B962B961B960B95FB95EB95DB95C",
		x"B97BB97AB979B978B977B976B975B974B973B972B971B970B96FB96EB96DB96C",
		x"B987B986B985B984B983B982B981B980FFFFFFFFFFFFFFFFB97FB97EB97DB97C",
		x"B997B996B995B994B993B992B991B990B98FB98EB98DB98CB98BB98AB989B988",
		x"B9A7B9A6B9A5B9A4B9A3B9A2B9A1B9A0B99FB99EB99DB99CB99BB99AB999B998",
		x"B9B7B9B6B9B5B9B4B9B3B9B2B9B1B9B0B9AFB9AEB9ADB9ACB9ABB9AAB9A9B9A8",
		x"B9C3B9C2B9C1B9C0FFFFFFFFFFFFFFFFB9BFB9BEB9BDB9BCB9BBB9BAB9B9B9B8",
		x"B9D3B9D2B9D1B9D0B9CFB9CEB9CDB9CCB9CBB9CAB9C9B9C8B9C7B9C6B9C5B9C4",
		x"B9E3B9E2B9E1B9E0B9DFB9DEB9DDB9DCB9DBB9DAB9D9B9D8B9D7B9D6B9D5B9D4",
		x"B9F3B9F2B9F1B9F0B9EFB9EEB9EDB9ECB9EBB9EAB9E9B9E8B9E7B9E6B9E5B9E4",
		x"FFFFFFFFFFFFFFFFB9FFB9FEB9FDB9FCB9FBB9FAB9F9B9F8B9F7B9F6B9F5B9F4",
		x"BA0FBA0EBA0DBA0CBA0BBA0ABA09BA08BA07BA06BA05BA04BA03BA02BA01BA00",
		x"BA1FBA1EBA1DBA1CBA1BBA1ABA19BA18BA17BA16BA15BA14BA13BA12BA11BA10",
		x"BA2FBA2EBA2DBA2CBA2BBA2ABA29BA28BA27BA26BA25BA24BA23BA22BA21BA20",
		x"BA3FBA3EBA3DBA3CBA3BBA3ABA39BA38BA37BA36BA35BA34BA33BA32BA31BA30",
		x"BA4BBA4ABA49BA48BA47BA46BA45BA44BA43BA42BA41BA40FFFFFFFFFFFFFFFF",
		x"BA5BBA5ABA59BA58BA57BA56BA55BA54BA53BA52BA51BA50BA4FBA4EBA4DBA4C",
		x"BA6BBA6ABA69BA68BA67BA66BA65BA64BA63BA62BA61BA60BA5FBA5EBA5DBA5C",
		x"BA7BBA7ABA79BA78BA77BA76BA75BA74BA73BA72BA71BA70BA6FBA6EBA6DBA6C",
		x"BA87BA86BA85BA84BA83BA82BA81BA80FFFFFFFFFFFFFFFFBA7FBA7EBA7DBA7C",
		x"BA97BA96BA95BA94BA93BA92BA91BA90BA8FBA8EBA8DBA8CBA8BBA8ABA89BA88",
		x"BAA7BAA6BAA5BAA4BAA3BAA2BAA1BAA0BA9FBA9EBA9DBA9CBA9BBA9ABA99BA98",
		x"BAB7BAB6BAB5BAB4BAB3BAB2BAB1BAB0BAAFBAAEBAADBAACBAABBAAABAA9BAA8",
		x"BAC3BAC2BAC1BAC0FFFFFFFFFFFFFFFFBABFBABEBABDBABCBABBBABABAB9BAB8",
		x"BAD3BAD2BAD1BAD0BACFBACEBACDBACCBACBBACABAC9BAC8BAC7BAC6BAC5BAC4",
		x"BAE3BAE2BAE1BAE0BADFBADEBADDBADCBADBBADABAD9BAD8BAD7BAD6BAD5BAD4",
		x"BAF3BAF2BAF1BAF0BAEFBAEEBAEDBAECBAEBBAEABAE9BAE8BAE7BAE6BAE5BAE4",
		x"FFFFFFFFFFFFFFFFBAFFBAFEBAFDBAFCBAFBBAFABAF9BAF8BAF7BAF6BAF5BAF4",
		x"BB0FBB0EBB0DBB0CBB0BBB0ABB09BB08BB07BB06BB05BB04BB03BB02BB01BB00",
		x"BB1FBB1EBB1DBB1CBB1BBB1ABB19BB18BB17BB16BB15BB14BB13BB12BB11BB10",
		x"BB2FBB2EBB2DBB2CBB2BBB2ABB29BB28BB27BB26BB25BB24BB23BB22BB21BB20",
		x"BB3FBB3EBB3DBB3CBB3BBB3ABB39BB38BB37BB36BB35BB34BB33BB32BB31BB30",
		x"BB4BBB4ABB49BB48BB47BB46BB45BB44BB43BB42BB41BB40FFFFFFFFFFFFFFFF",
		x"BB5BBB5ABB59BB58BB57BB56BB55BB54BB53BB52BB51BB50BB4FBB4EBB4DBB4C",
		x"BB6BBB6ABB69BB68BB67BB66BB65BB64BB63BB62BB61BB60BB5FBB5EBB5DBB5C",
		x"BB7BBB7ABB79BB78BB77BB76BB75BB74BB73BB72BB71BB70BB6FBB6EBB6DBB6C",
		x"BB87BB86BB85BB84BB83BB82BB81BB80FFFFFFFFFFFFFFFFBB7FBB7EBB7DBB7C",
		x"BB97BB96BB95BB94BB93BB92BB91BB90BB8FBB8EBB8DBB8CBB8BBB8ABB89BB88",
		x"BBA7BBA6BBA5BBA4BBA3BBA2BBA1BBA0BB9FBB9EBB9DBB9CBB9BBB9ABB99BB98",
		x"BBB7BBB6BBB5BBB4BBB3BBB2BBB1BBB0BBAFBBAEBBADBBACBBABBBAABBA9BBA8",
		x"BBC3BBC2BBC1BBC0FFFFFFFFFFFFFFFFBBBFBBBEBBBDBBBCBBBBBBBABBB9BBB8",
		x"BBD3BBD2BBD1BBD0BBCFBBCEBBCDBBCCBBCBBBCABBC9BBC8BBC7BBC6BBC5BBC4",
		x"BBE3BBE2BBE1BBE0BBDFBBDEBBDDBBDCBBDBBBDABBD9BBD8BBD7BBD6BBD5BBD4",
		x"BBF3BBF2BBF1BBF0BBEFBBEEBBEDBBECBBEBBBEABBE9BBE8BBE7BBE6BBE5BBE4",
		x"FFFFFFFFFFFFFFFFBBFFBBFEBBFDBBFCBBFBBBFABBF9BBF8BBF7BBF6BBF5BBF4",
		x"BC0FBC0EBC0DBC0CBC0BBC0ABC09BC08BC07BC06BC05BC04BC03BC02BC01BC00",
		x"BC1FBC1EBC1DBC1CBC1BBC1ABC19BC18BC17BC16BC15BC14BC13BC12BC11BC10",
		x"BC2FBC2EBC2DBC2CBC2BBC2ABC29BC28BC27BC26BC25BC24BC23BC22BC21BC20",
		x"BC3FBC3EBC3DBC3CBC3BBC3ABC39BC38BC37BC36BC35BC34BC33BC32BC31BC30",
		x"BC4BBC4ABC49BC48BC47BC46BC45BC44BC43BC42BC41BC40FFFFFFFFFFFFFFFF",
		x"BC5BBC5ABC59BC58BC57BC56BC55BC54BC53BC52BC51BC50BC4FBC4EBC4DBC4C",
		x"BC6BBC6ABC69BC68BC67BC66BC65BC64BC63BC62BC61BC60BC5FBC5EBC5DBC5C",
		x"BC7BBC7ABC79BC78BC77BC76BC75BC74BC73BC72BC71BC70BC6FBC6EBC6DBC6C",
		x"BC87BC86BC85BC84BC83BC82BC81BC80FFFFFFFFFFFFFFFFBC7FBC7EBC7DBC7C",
		x"BC97BC96BC95BC94BC93BC92BC91BC90BC8FBC8EBC8DBC8CBC8BBC8ABC89BC88",
		x"BCA7BCA6BCA5BCA4BCA3BCA2BCA1BCA0BC9FBC9EBC9DBC9CBC9BBC9ABC99BC98",
		x"BCB7BCB6BCB5BCB4BCB3BCB2BCB1BCB0BCAFBCAEBCADBCACBCABBCAABCA9BCA8",
		x"BCC3BCC2BCC1BCC0FFFFFFFFFFFFFFFFBCBFBCBEBCBDBCBCBCBBBCBABCB9BCB8",
		x"BCD3BCD2BCD1BCD0BCCFBCCEBCCDBCCCBCCBBCCABCC9BCC8BCC7BCC6BCC5BCC4",
		x"BCE3BCE2BCE1BCE0BCDFBCDEBCDDBCDCBCDBBCDABCD9BCD8BCD7BCD6BCD5BCD4",
		x"BCF3BCF2BCF1BCF0BCEFBCEEBCEDBCECBCEBBCEABCE9BCE8BCE7BCE6BCE5BCE4",
		x"FFFFFFFFFFFFFFFFBCFFBCFEBCFDBCFCBCFBBCFABCF9BCF8BCF7BCF6BCF5BCF4",
		x"BD0FBD0EBD0DBD0CBD0BBD0ABD09BD08BD07BD06BD05BD04BD03BD02BD01BD00",
		x"BD1FBD1EBD1DBD1CBD1BBD1ABD19BD18BD17BD16BD15BD14BD13BD12BD11BD10",
		x"BD2FBD2EBD2DBD2CBD2BBD2ABD29BD28BD27BD26BD25BD24BD23BD22BD21BD20",
		x"BD3FBD3EBD3DBD3CBD3BBD3ABD39BD38BD37BD36BD35BD34BD33BD32BD31BD30",
		x"BD4BBD4ABD49BD48BD47BD46BD45BD44BD43BD42BD41BD40FFFFFFFFFFFFFFFF",
		x"BD5BBD5ABD59BD58BD57BD56BD55BD54BD53BD52BD51BD50BD4FBD4EBD4DBD4C",
		x"BD6BBD6ABD69BD68BD67BD66BD65BD64BD63BD62BD61BD60BD5FBD5EBD5DBD5C",
		x"BD7BBD7ABD79BD78BD77BD76BD75BD74BD73BD72BD71BD70BD6FBD6EBD6DBD6C",
		x"BD87BD86BD85BD84BD83BD82BD81BD80FFFFFFFFFFFFFFFFBD7FBD7EBD7DBD7C",
		x"BD97BD96BD95BD94BD93BD92BD91BD90BD8FBD8EBD8DBD8CBD8BBD8ABD89BD88",
		x"BDA7BDA6BDA5BDA4BDA3BDA2BDA1BDA0BD9FBD9EBD9DBD9CBD9BBD9ABD99BD98",
		x"BDB7BDB6BDB5BDB4BDB3BDB2BDB1BDB0BDAFBDAEBDADBDACBDABBDAABDA9BDA8",
		x"BDC3BDC2BDC1BDC0FFFFFFFFFFFFFFFFBDBFBDBEBDBDBDBCBDBBBDBABDB9BDB8",
		x"BDD3BDD2BDD1BDD0BDCFBDCEBDCDBDCCBDCBBDCABDC9BDC8BDC7BDC6BDC5BDC4",
		x"BDE3BDE2BDE1BDE0BDDFBDDEBDDDBDDCBDDBBDDABDD9BDD8BDD7BDD6BDD5BDD4",
		x"BDF3BDF2BDF1BDF0BDEFBDEEBDEDBDECBDEBBDEABDE9BDE8BDE7BDE6BDE5BDE4",
		x"FFFFFFFFFFFFFFFFBDFFBDFEBDFDBDFCBDFBBDFABDF9BDF8BDF7BDF6BDF5BDF4",
		x"BE0FBE0EBE0DBE0CBE0BBE0ABE09BE08BE07BE06BE05BE04BE03BE02BE01BE00",
		x"BE1FBE1EBE1DBE1CBE1BBE1ABE19BE18BE17BE16BE15BE14BE13BE12BE11BE10",
		x"BE2FBE2EBE2DBE2CBE2BBE2ABE29BE28BE27BE26BE25BE24BE23BE22BE21BE20",
		x"BE3FBE3EBE3DBE3CBE3BBE3ABE39BE38BE37BE36BE35BE34BE33BE32BE31BE30",
		x"BE4BBE4ABE49BE48BE47BE46BE45BE44BE43BE42BE41BE40FFFFFFFFFFFFFFFF",
		x"BE5BBE5ABE59BE58BE57BE56BE55BE54BE53BE52BE51BE50BE4FBE4EBE4DBE4C",
		x"BE6BBE6ABE69BE68BE67BE66BE65BE64BE63BE62BE61BE60BE5FBE5EBE5DBE5C",
		x"BE7BBE7ABE79BE78BE77BE76BE75BE74BE73BE72BE71BE70BE6FBE6EBE6DBE6C",
		x"BE87BE86BE85BE84BE83BE82BE81BE80FFFFFFFFFFFFFFFFBE7FBE7EBE7DBE7C",
		x"BE97BE96BE95BE94BE93BE92BE91BE90BE8FBE8EBE8DBE8CBE8BBE8ABE89BE88",
		x"BEA7BEA6BEA5BEA4BEA3BEA2BEA1BEA0BE9FBE9EBE9DBE9CBE9BBE9ABE99BE98",
		x"BEB7BEB6BEB5BEB4BEB3BEB2BEB1BEB0BEAFBEAEBEADBEACBEABBEAABEA9BEA8",
		x"BEC3BEC2BEC1BEC0FFFFFFFFFFFFFFFFBEBFBEBEBEBDBEBCBEBBBEBABEB9BEB8",
		x"BED3BED2BED1BED0BECFBECEBECDBECCBECBBECABEC9BEC8BEC7BEC6BEC5BEC4",
		x"BEE3BEE2BEE1BEE0BEDFBEDEBEDDBEDCBEDBBEDABED9BED8BED7BED6BED5BED4",
		x"BEF3BEF2BEF1BEF0BEEFBEEEBEEDBEECBEEBBEEABEE9BEE8BEE7BEE6BEE5BEE4",
		x"FFFFFFFFFFFFFFFFBEFFBEFEBEFDBEFCBEFBBEFABEF9BEF8BEF7BEF6BEF5BEF4",
		x"BF0FBF0EBF0DBF0CBF0BBF0ABF09BF08BF07BF06BF05BF04BF03BF02BF01BF00",
		x"BF1FBF1EBF1DBF1CBF1BBF1ABF19BF18BF17BF16BF15BF14BF13BF12BF11BF10",
		x"BF2FBF2EBF2DBF2CBF2BBF2ABF29BF28BF27BF26BF25BF24BF23BF22BF21BF20",
		x"BF3FBF3EBF3DBF3CBF3BBF3ABF39BF38BF37BF36BF35BF34BF33BF32BF31BF30",
		x"BF4BBF4ABF49BF48BF47BF46BF45BF44BF43BF42BF41BF40FFFFFFFFFFFFFFFF",
		x"BF5BBF5ABF59BF58BF57BF56BF55BF54BF53BF52BF51BF50BF4FBF4EBF4DBF4C",
		x"BF6BBF6ABF69BF68BF67BF66BF65BF64BF63BF62BF61BF60BF5FBF5EBF5DBF5C",
		x"BF7BBF7ABF79BF78BF77BF76BF75BF74BF73BF72BF71BF70BF6FBF6EBF6DBF6C",
		x"BF87BF86BF85BF84BF83BF82BF81BF80FFFFFFFFFFFFFFFFBF7FBF7EBF7DBF7C",
		x"BF97BF96BF95BF94BF93BF92BF91BF90BF8FBF8EBF8DBF8CBF8BBF8ABF89BF88",
		x"BFA7BFA6BFA5BFA4BFA3BFA2BFA1BFA0BF9FBF9EBF9DBF9CBF9BBF9ABF99BF98",
		x"BFB7BFB6BFB5BFB4BFB3BFB2BFB1BFB0BFAFBFAEBFADBFACBFABBFAABFA9BFA8",
		x"BFC3BFC2BFC1BFC0FFFFFFFFFFFFFFFFBFBFBFBEBFBDBFBCBFBBBFBABFB9BFB8",
		x"BFD3BFD2BFD1BFD0BFCFBFCEBFCDBFCCBFCBBFCABFC9BFC8BFC7BFC6BFC5BFC4",
		x"BFE3BFE2BFE1BFE0BFDFBFDEBFDDBFDCBFDBBFDABFD9BFD8BFD7BFD6BFD5BFD4",
		x"BFF3BFF2BFF1BFF0BFEFBFEEBFEDBFECBFEBBFEABFE9BFE8BFE7BFE6BFE5BFE4",
		x"FFFFFFFFFFFFFFFFBFFFBFFEBFFDBFFCBFFBBFFABFF9BFF8BFF7BFF6BFF5BFF4",
		x"C00FC00EC00DC00CC00BC00AC009C008C007C006C005C004C003C002C001C000",
		x"C01FC01EC01DC01CC01BC01AC019C018C017C016C015C014C013C012C011C010",
		x"C02FC02EC02DC02CC02BC02AC029C028C027C026C025C024C023C022C021C020",
		x"C03FC03EC03DC03CC03BC03AC039C038C037C036C035C034C033C032C031C030",
		x"C04BC04AC049C048C047C046C045C044C043C042C041C040FFFFFFFFFFFFFFFF",
		x"C05BC05AC059C058C057C056C055C054C053C052C051C050C04FC04EC04DC04C",
		x"C06BC06AC069C068C067C066C065C064C063C062C061C060C05FC05EC05DC05C",
		x"C07BC07AC079C078C077C076C075C074C073C072C071C070C06FC06EC06DC06C",
		x"C087C086C085C084C083C082C081C080FFFFFFFFFFFFFFFFC07FC07EC07DC07C",
		x"C097C096C095C094C093C092C091C090C08FC08EC08DC08CC08BC08AC089C088",
		x"C0A7C0A6C0A5C0A4C0A3C0A2C0A1C0A0C09FC09EC09DC09CC09BC09AC099C098",
		x"C0B7C0B6C0B5C0B4C0B3C0B2C0B1C0B0C0AFC0AEC0ADC0ACC0ABC0AAC0A9C0A8",
		x"C0C3C0C2C0C1C0C0FFFFFFFFFFFFFFFFC0BFC0BEC0BDC0BCC0BBC0BAC0B9C0B8",
		x"C0D3C0D2C0D1C0D0C0CFC0CEC0CDC0CCC0CBC0CAC0C9C0C8C0C7C0C6C0C5C0C4",
		x"C0E3C0E2C0E1C0E0C0DFC0DEC0DDC0DCC0DBC0DAC0D9C0D8C0D7C0D6C0D5C0D4",
		x"C0F3C0F2C0F1C0F0C0EFC0EEC0EDC0ECC0EBC0EAC0E9C0E8C0E7C0E6C0E5C0E4",
		x"FFFFFFFFFFFFFFFFC0FFC0FEC0FDC0FCC0FBC0FAC0F9C0F8C0F7C0F6C0F5C0F4",
		x"C10FC10EC10DC10CC10BC10AC109C108C107C106C105C104C103C102C101C100",
		x"C11FC11EC11DC11CC11BC11AC119C118C117C116C115C114C113C112C111C110",
		x"C12FC12EC12DC12CC12BC12AC129C128C127C126C125C124C123C122C121C120",
		x"C13FC13EC13DC13CC13BC13AC139C138C137C136C135C134C133C132C131C130",
		x"C14BC14AC149C148C147C146C145C144C143C142C141C140FFFFFFFFFFFFFFFF",
		x"C15BC15AC159C158C157C156C155C154C153C152C151C150C14FC14EC14DC14C",
		x"C16BC16AC169C168C167C166C165C164C163C162C161C160C15FC15EC15DC15C",
		x"C17BC17AC179C178C177C176C175C174C173C172C171C170C16FC16EC16DC16C",
		x"C187C186C185C184C183C182C181C180FFFFFFFFFFFFFFFFC17FC17EC17DC17C",
		x"C197C196C195C194C193C192C191C190C18FC18EC18DC18CC18BC18AC189C188",
		x"C1A7C1A6C1A5C1A4C1A3C1A2C1A1C1A0C19FC19EC19DC19CC19BC19AC199C198",
		x"C1B7C1B6C1B5C1B4C1B3C1B2C1B1C1B0C1AFC1AEC1ADC1ACC1ABC1AAC1A9C1A8",
		x"C1C3C1C2C1C1C1C0FFFFFFFFFFFFFFFFC1BFC1BEC1BDC1BCC1BBC1BAC1B9C1B8",
		x"C1D3C1D2C1D1C1D0C1CFC1CEC1CDC1CCC1CBC1CAC1C9C1C8C1C7C1C6C1C5C1C4",
		x"C1E3C1E2C1E1C1E0C1DFC1DEC1DDC1DCC1DBC1DAC1D9C1D8C1D7C1D6C1D5C1D4",
		x"C1F3C1F2C1F1C1F0C1EFC1EEC1EDC1ECC1EBC1EAC1E9C1E8C1E7C1E6C1E5C1E4",
		x"FFFFFFFFFFFFFFFFC1FFC1FEC1FDC1FCC1FBC1FAC1F9C1F8C1F7C1F6C1F5C1F4",
		x"C20FC20EC20DC20CC20BC20AC209C208C207C206C205C204C203C202C201C200",
		x"C21FC21EC21DC21CC21BC21AC219C218C217C216C215C214C213C212C211C210",
		x"C22FC22EC22DC22CC22BC22AC229C228C227C226C225C224C223C222C221C220",
		x"C23FC23EC23DC23CC23BC23AC239C238C237C236C235C234C233C232C231C230",
		x"C24BC24AC249C248C247C246C245C244C243C242C241C240FFFFFFFFFFFFFFFF",
		x"C25BC25AC259C258C257C256C255C254C253C252C251C250C24FC24EC24DC24C",
		x"C26BC26AC269C268C267C266C265C264C263C262C261C260C25FC25EC25DC25C",
		x"C27BC27AC279C278C277C276C275C274C273C272C271C270C26FC26EC26DC26C",
		x"C287C286C285C284C283C282C281C280FFFFFFFFFFFFFFFFC27FC27EC27DC27C",
		x"C297C296C295C294C293C292C291C290C28FC28EC28DC28CC28BC28AC289C288",
		x"C2A7C2A6C2A5C2A4C2A3C2A2C2A1C2A0C29FC29EC29DC29CC29BC29AC299C298",
		x"C2B7C2B6C2B5C2B4C2B3C2B2C2B1C2B0C2AFC2AEC2ADC2ACC2ABC2AAC2A9C2A8",
		x"C2C3C2C2C2C1C2C0FFFFFFFFFFFFFFFFC2BFC2BEC2BDC2BCC2BBC2BAC2B9C2B8",
		x"C2D3C2D2C2D1C2D0C2CFC2CEC2CDC2CCC2CBC2CAC2C9C2C8C2C7C2C6C2C5C2C4",
		x"C2E3C2E2C2E1C2E0C2DFC2DEC2DDC2DCC2DBC2DAC2D9C2D8C2D7C2D6C2D5C2D4",
		x"C2F3C2F2C2F1C2F0C2EFC2EEC2EDC2ECC2EBC2EAC2E9C2E8C2E7C2E6C2E5C2E4",
		x"FFFFFFFFFFFFFFFFC2FFC2FEC2FDC2FCC2FBC2FAC2F9C2F8C2F7C2F6C2F5C2F4",
		x"C30FC30EC30DC30CC30BC30AC309C308C307C306C305C304C303C302C301C300",
		x"C31FC31EC31DC31CC31BC31AC319C318C317C316C315C314C313C312C311C310",
		x"C32FC32EC32DC32CC32BC32AC329C328C327C326C325C324C323C322C321C320",
		x"C33FC33EC33DC33CC33BC33AC339C338C337C336C335C334C333C332C331C330",
		x"C34BC34AC349C348C347C346C345C344C343C342C341C340FFFFFFFFFFFFFFFF",
		x"C35BC35AC359C358C357C356C355C354C353C352C351C350C34FC34EC34DC34C",
		x"C36BC36AC369C368C367C366C365C364C363C362C361C360C35FC35EC35DC35C",
		x"C37BC37AC379C378C377C376C375C374C373C372C371C370C36FC36EC36DC36C",
		x"C387C386C385C384C383C382C381C380FFFFFFFFFFFFFFFFC37FC37EC37DC37C",
		x"C397C396C395C394C393C392C391C390C38FC38EC38DC38CC38BC38AC389C388",
		x"C3A7C3A6C3A5C3A4C3A3C3A2C3A1C3A0C39FC39EC39DC39CC39BC39AC399C398",
		x"C3B7C3B6C3B5C3B4C3B3C3B2C3B1C3B0C3AFC3AEC3ADC3ACC3ABC3AAC3A9C3A8",
		x"C3C3C3C2C3C1C3C0FFFFFFFFFFFFFFFFC3BFC3BEC3BDC3BCC3BBC3BAC3B9C3B8",
		x"C3D3C3D2C3D1C3D0C3CFC3CEC3CDC3CCC3CBC3CAC3C9C3C8C3C7C3C6C3C5C3C4",
		x"C3E3C3E2C3E1C3E0C3DFC3DEC3DDC3DCC3DBC3DAC3D9C3D8C3D7C3D6C3D5C3D4",
		x"C3F3C3F2C3F1C3F0C3EFC3EEC3EDC3ECC3EBC3EAC3E9C3E8C3E7C3E6C3E5C3E4",
		x"FFFFFFFFFFFFFFFFC3FFC3FEC3FDC3FCC3FBC3FAC3F9C3F8C3F7C3F6C3F5C3F4",
		x"C40FC40EC40DC40CC40BC40AC409C408C407C406C405C404C403C402C401C400",
		x"C41FC41EC41DC41CC41BC41AC419C418C417C416C415C414C413C412C411C410",
		x"C42FC42EC42DC42CC42BC42AC429C428C427C426C425C424C423C422C421C420",
		x"C43FC43EC43DC43CC43BC43AC439C438C437C436C435C434C433C432C431C430",
		x"C44BC44AC449C448C447C446C445C444C443C442C441C440FFFFFFFFFFFFFFFF",
		x"C45BC45AC459C458C457C456C455C454C453C452C451C450C44FC44EC44DC44C",
		x"C46BC46AC469C468C467C466C465C464C463C462C461C460C45FC45EC45DC45C",
		x"C47BC47AC479C478C477C476C475C474C473C472C471C470C46FC46EC46DC46C",
		x"C487C486C485C484C483C482C481C480FFFFFFFFFFFFFFFFC47FC47EC47DC47C",
		x"C497C496C495C494C493C492C491C490C48FC48EC48DC48CC48BC48AC489C488",
		x"C4A7C4A6C4A5C4A4C4A3C4A2C4A1C4A0C49FC49EC49DC49CC49BC49AC499C498",
		x"C4B7C4B6C4B5C4B4C4B3C4B2C4B1C4B0C4AFC4AEC4ADC4ACC4ABC4AAC4A9C4A8",
		x"C4C3C4C2C4C1C4C0FFFFFFFFFFFFFFFFC4BFC4BEC4BDC4BCC4BBC4BAC4B9C4B8",
		x"C4D3C4D2C4D1C4D0C4CFC4CEC4CDC4CCC4CBC4CAC4C9C4C8C4C7C4C6C4C5C4C4",
		x"C4E3C4E2C4E1C4E0C4DFC4DEC4DDC4DCC4DBC4DAC4D9C4D8C4D7C4D6C4D5C4D4",
		x"C4F3C4F2C4F1C4F0C4EFC4EEC4EDC4ECC4EBC4EAC4E9C4E8C4E7C4E6C4E5C4E4",
		x"FFFFFFFFFFFFFFFFC4FFC4FEC4FDC4FCC4FBC4FAC4F9C4F8C4F7C4F6C4F5C4F4",
		x"C50FC50EC50DC50CC50BC50AC509C508C507C506C505C504C503C502C501C500",
		x"C51FC51EC51DC51CC51BC51AC519C518C517C516C515C514C513C512C511C510",
		x"C52FC52EC52DC52CC52BC52AC529C528C527C526C525C524C523C522C521C520",
		x"C53FC53EC53DC53CC53BC53AC539C538C537C536C535C534C533C532C531C530",
		x"C54BC54AC549C548C547C546C545C544C543C542C541C540FFFFFFFFFFFFFFFF",
		x"C55BC55AC559C558C557C556C555C554C553C552C551C550C54FC54EC54DC54C",
		x"C56BC56AC569C568C567C566C565C564C563C562C561C560C55FC55EC55DC55C",
		x"C57BC57AC579C578C577C576C575C574C573C572C571C570C56FC56EC56DC56C",
		x"C587C586C585C584C583C582C581C580FFFFFFFFFFFFFFFFC57FC57EC57DC57C",
		x"C597C596C595C594C593C592C591C590C58FC58EC58DC58CC58BC58AC589C588",
		x"C5A7C5A6C5A5C5A4C5A3C5A2C5A1C5A0C59FC59EC59DC59CC59BC59AC599C598",
		x"C5B7C5B6C5B5C5B4C5B3C5B2C5B1C5B0C5AFC5AEC5ADC5ACC5ABC5AAC5A9C5A8",
		x"C5C3C5C2C5C1C5C0FFFFFFFFFFFFFFFFC5BFC5BEC5BDC5BCC5BBC5BAC5B9C5B8",
		x"C5D3C5D2C5D1C5D0C5CFC5CEC5CDC5CCC5CBC5CAC5C9C5C8C5C7C5C6C5C5C5C4",
		x"C5E3C5E2C5E1C5E0C5DFC5DEC5DDC5DCC5DBC5DAC5D9C5D8C5D7C5D6C5D5C5D4",
		x"C5F3C5F2C5F1C5F0C5EFC5EEC5EDC5ECC5EBC5EAC5E9C5E8C5E7C5E6C5E5C5E4",
		x"FFFFFFFFFFFFFFFFC5FFC5FEC5FDC5FCC5FBC5FAC5F9C5F8C5F7C5F6C5F5C5F4",
		x"C60FC60EC60DC60CC60BC60AC609C608C607C606C605C604C603C602C601C600",
		x"C61FC61EC61DC61CC61BC61AC619C618C617C616C615C614C613C612C611C610",
		x"C62FC62EC62DC62CC62BC62AC629C628C627C626C625C624C623C622C621C620",
		x"C63FC63EC63DC63CC63BC63AC639C638C637C636C635C634C633C632C631C630",
		x"C64BC64AC649C648C647C646C645C644C643C642C641C640FFFFFFFFFFFFFFFF",
		x"C65BC65AC659C658C657C656C655C654C653C652C651C650C64FC64EC64DC64C",
		x"C66BC66AC669C668C667C666C665C664C663C662C661C660C65FC65EC65DC65C",
		x"C67BC67AC679C678C677C676C675C674C673C672C671C670C66FC66EC66DC66C",
		x"C687C686C685C684C683C682C681C680FFFFFFFFFFFFFFFFC67FC67EC67DC67C",
		x"C697C696C695C694C693C692C691C690C68FC68EC68DC68CC68BC68AC689C688",
		x"C6A7C6A6C6A5C6A4C6A3C6A2C6A1C6A0C69FC69EC69DC69CC69BC69AC699C698",
		x"C6B7C6B6C6B5C6B4C6B3C6B2C6B1C6B0C6AFC6AEC6ADC6ACC6ABC6AAC6A9C6A8",
		x"C6C3C6C2C6C1C6C0FFFFFFFFFFFFFFFFC6BFC6BEC6BDC6BCC6BBC6BAC6B9C6B8",
		x"C6D3C6D2C6D1C6D0C6CFC6CEC6CDC6CCC6CBC6CAC6C9C6C8C6C7C6C6C6C5C6C4",
		x"C6E3C6E2C6E1C6E0C6DFC6DEC6DDC6DCC6DBC6DAC6D9C6D8C6D7C6D6C6D5C6D4",
		x"C6F3C6F2C6F1C6F0C6EFC6EEC6EDC6ECC6EBC6EAC6E9C6E8C6E7C6E6C6E5C6E4",
		x"FFFFFFFFFFFFFFFFC6FFC6FEC6FDC6FCC6FBC6FAC6F9C6F8C6F7C6F6C6F5C6F4",
		x"C70FC70EC70DC70CC70BC70AC709C708C707C706C705C704C703C702C701C700",
		x"C71FC71EC71DC71CC71BC71AC719C718C717C716C715C714C713C712C711C710",
		x"C72FC72EC72DC72CC72BC72AC729C728C727C726C725C724C723C722C721C720",
		x"C73FC73EC73DC73CC73BC73AC739C738C737C736C735C734C733C732C731C730",
		x"C74BC74AC749C748C747C746C745C744C743C742C741C740FFFFFFFFFFFFFFFF",
		x"C75BC75AC759C758C757C756C755C754C753C752C751C750C74FC74EC74DC74C",
		x"C76BC76AC769C768C767C766C765C764C763C762C761C760C75FC75EC75DC75C",
		x"C77BC77AC779C778C777C776C775C774C773C772C771C770C76FC76EC76DC76C",
		x"C787C786C785C784C783C782C781C780FFFFFFFFFFFFFFFFC77FC77EC77DC77C",
		x"C797C796C795C794C793C792C791C790C78FC78EC78DC78CC78BC78AC789C788",
		x"C7A7C7A6C7A5C7A4C7A3C7A2C7A1C7A0C79FC79EC79DC79CC79BC79AC799C798",
		x"C7B7C7B6C7B5C7B4C7B3C7B2C7B1C7B0C7AFC7AEC7ADC7ACC7ABC7AAC7A9C7A8",
		x"C7C3C7C2C7C1C7C0FFFFFFFFFFFFFFFFC7BFC7BEC7BDC7BCC7BBC7BAC7B9C7B8",
		x"C7D3C7D2C7D1C7D0C7CFC7CEC7CDC7CCC7CBC7CAC7C9C7C8C7C7C7C6C7C5C7C4",
		x"C7E3C7E2C7E1C7E0C7DFC7DEC7DDC7DCC7DBC7DAC7D9C7D8C7D7C7D6C7D5C7D4",
		x"C7F3C7F2C7F1C7F0C7EFC7EEC7EDC7ECC7EBC7EAC7E9C7E8C7E7C7E6C7E5C7E4",
		x"FFFFFFFFFFFFFFFFC7FFC7FEC7FDC7FCC7FBC7FAC7F9C7F8C7F7C7F6C7F5C7F4",
		x"C80FC80EC80DC80CC80BC80AC809C808C807C806C805C804C803C802C801C800",
		x"C81FC81EC81DC81CC81BC81AC819C818C817C816C815C814C813C812C811C810",
		x"C82FC82EC82DC82CC82BC82AC829C828C827C826C825C824C823C822C821C820",
		x"C83FC83EC83DC83CC83BC83AC839C838C837C836C835C834C833C832C831C830",
		x"C84BC84AC849C848C847C846C845C844C843C842C841C840FFFFFFFFFFFFFFFF",
		x"C85BC85AC859C858C857C856C855C854C853C852C851C850C84FC84EC84DC84C",
		x"C86BC86AC869C868C867C866C865C864C863C862C861C860C85FC85EC85DC85C",
		x"C87BC87AC879C878C877C876C875C874C873C872C871C870C86FC86EC86DC86C",
		x"C887C886C885C884C883C882C881C880FFFFFFFFFFFFFFFFC87FC87EC87DC87C",
		x"C897C896C895C894C893C892C891C890C88FC88EC88DC88CC88BC88AC889C888",
		x"C8A7C8A6C8A5C8A4C8A3C8A2C8A1C8A0C89FC89EC89DC89CC89BC89AC899C898",
		x"C8B7C8B6C8B5C8B4C8B3C8B2C8B1C8B0C8AFC8AEC8ADC8ACC8ABC8AAC8A9C8A8",
		x"C8C3C8C2C8C1C8C0FFFFFFFFFFFFFFFFC8BFC8BEC8BDC8BCC8BBC8BAC8B9C8B8",
		x"C8D3C8D2C8D1C8D0C8CFC8CEC8CDC8CCC8CBC8CAC8C9C8C8C8C7C8C6C8C5C8C4",
		x"C8E3C8E2C8E1C8E0C8DFC8DEC8DDC8DCC8DBC8DAC8D9C8D8C8D7C8D6C8D5C8D4",
		x"C8F3C8F2C8F1C8F0C8EFC8EEC8EDC8ECC8EBC8EAC8E9C8E8C8E7C8E6C8E5C8E4",
		x"FFFFFFFFFFFFFFFFC8FFC8FEC8FDC8FCC8FBC8FAC8F9C8F8C8F7C8F6C8F5C8F4",
		x"C90FC90EC90DC90CC90BC90AC909C908C907C906C905C904C903C902C901C900",
		x"C91FC91EC91DC91CC91BC91AC919C918C917C916C915C914C913C912C911C910",
		x"C92FC92EC92DC92CC92BC92AC929C928C927C926C925C924C923C922C921C920",
		x"C93FC93EC93DC93CC93BC93AC939C938C937C936C935C934C933C932C931C930",
		x"C94BC94AC949C948C947C946C945C944C943C942C941C940FFFFFFFFFFFFFFFF",
		x"C95BC95AC959C958C957C956C955C954C953C952C951C950C94FC94EC94DC94C",
		x"C96BC96AC969C968C967C966C965C964C963C962C961C960C95FC95EC95DC95C",
		x"C97BC97AC979C978C977C976C975C974C973C972C971C970C96FC96EC96DC96C",
		x"C987C986C985C984C983C982C981C980FFFFFFFFFFFFFFFFC97FC97EC97DC97C",
		x"C997C996C995C994C993C992C991C990C98FC98EC98DC98CC98BC98AC989C988",
		x"C9A7C9A6C9A5C9A4C9A3C9A2C9A1C9A0C99FC99EC99DC99CC99BC99AC999C998",
		x"C9B7C9B6C9B5C9B4C9B3C9B2C9B1C9B0C9AFC9AEC9ADC9ACC9ABC9AAC9A9C9A8",
		x"C9C3C9C2C9C1C9C0FFFFFFFFFFFFFFFFC9BFC9BEC9BDC9BCC9BBC9BAC9B9C9B8",
		x"C9D3C9D2C9D1C9D0C9CFC9CEC9CDC9CCC9CBC9CAC9C9C9C8C9C7C9C6C9C5C9C4",
		x"C9E3C9E2C9E1C9E0C9DFC9DEC9DDC9DCC9DBC9DAC9D9C9D8C9D7C9D6C9D5C9D4",
		x"C9F3C9F2C9F1C9F0C9EFC9EEC9EDC9ECC9EBC9EAC9E9C9E8C9E7C9E6C9E5C9E4",
		x"FFFFFFFFFFFFFFFFC9FFC9FEC9FDC9FCC9FBC9FAC9F9C9F8C9F7C9F6C9F5C9F4",
		x"CA0FCA0ECA0DCA0CCA0BCA0ACA09CA08CA07CA06CA05CA04CA03CA02CA01CA00",
		x"CA1FCA1ECA1DCA1CCA1BCA1ACA19CA18CA17CA16CA15CA14CA13CA12CA11CA10",
		x"CA2FCA2ECA2DCA2CCA2BCA2ACA29CA28CA27CA26CA25CA24CA23CA22CA21CA20",
		x"CA3FCA3ECA3DCA3CCA3BCA3ACA39CA38CA37CA36CA35CA34CA33CA32CA31CA30",
		x"CA4BCA4ACA49CA48CA47CA46CA45CA44CA43CA42CA41CA40FFFFFFFFFFFFFFFF",
		x"CA5BCA5ACA59CA58CA57CA56CA55CA54CA53CA52CA51CA50CA4FCA4ECA4DCA4C",
		x"CA6BCA6ACA69CA68CA67CA66CA65CA64CA63CA62CA61CA60CA5FCA5ECA5DCA5C",
		x"CA7BCA7ACA79CA78CA77CA76CA75CA74CA73CA72CA71CA70CA6FCA6ECA6DCA6C",
		x"CA87CA86CA85CA84CA83CA82CA81CA80FFFFFFFFFFFFFFFFCA7FCA7ECA7DCA7C",
		x"CA97CA96CA95CA94CA93CA92CA91CA90CA8FCA8ECA8DCA8CCA8BCA8ACA89CA88",
		x"CAA7CAA6CAA5CAA4CAA3CAA2CAA1CAA0CA9FCA9ECA9DCA9CCA9BCA9ACA99CA98",
		x"CAB7CAB6CAB5CAB4CAB3CAB2CAB1CAB0CAAFCAAECAADCAACCAABCAAACAA9CAA8",
		x"CAC3CAC2CAC1CAC0FFFFFFFFFFFFFFFFCABFCABECABDCABCCABBCABACAB9CAB8",
		x"CAD3CAD2CAD1CAD0CACFCACECACDCACCCACBCACACAC9CAC8CAC7CAC6CAC5CAC4",
		x"CAE3CAE2CAE1CAE0CADFCADECADDCADCCADBCADACAD9CAD8CAD7CAD6CAD5CAD4",
		x"CAF3CAF2CAF1CAF0CAEFCAEECAEDCAECCAEBCAEACAE9CAE8CAE7CAE6CAE5CAE4",
		x"FFFFFFFFFFFFFFFFCAFFCAFECAFDCAFCCAFBCAFACAF9CAF8CAF7CAF6CAF5CAF4",
		x"CB0FCB0ECB0DCB0CCB0BCB0ACB09CB08CB07CB06CB05CB04CB03CB02CB01CB00",
		x"CB1FCB1ECB1DCB1CCB1BCB1ACB19CB18CB17CB16CB15CB14CB13CB12CB11CB10",
		x"CB2FCB2ECB2DCB2CCB2BCB2ACB29CB28CB27CB26CB25CB24CB23CB22CB21CB20",
		x"CB3FCB3ECB3DCB3CCB3BCB3ACB39CB38CB37CB36CB35CB34CB33CB32CB31CB30",
		x"CB4BCB4ACB49CB48CB47CB46CB45CB44CB43CB42CB41CB40FFFFFFFFFFFFFFFF",
		x"CB5BCB5ACB59CB58CB57CB56CB55CB54CB53CB52CB51CB50CB4FCB4ECB4DCB4C",
		x"CB6BCB6ACB69CB68CB67CB66CB65CB64CB63CB62CB61CB60CB5FCB5ECB5DCB5C",
		x"CB7BCB7ACB79CB78CB77CB76CB75CB74CB73CB72CB71CB70CB6FCB6ECB6DCB6C",
		x"CB87CB86CB85CB84CB83CB82CB81CB80FFFFFFFFFFFFFFFFCB7FCB7ECB7DCB7C",
		x"CB97CB96CB95CB94CB93CB92CB91CB90CB8FCB8ECB8DCB8CCB8BCB8ACB89CB88",
		x"CBA7CBA6CBA5CBA4CBA3CBA2CBA1CBA0CB9FCB9ECB9DCB9CCB9BCB9ACB99CB98",
		x"CBB7CBB6CBB5CBB4CBB3CBB2CBB1CBB0CBAFCBAECBADCBACCBABCBAACBA9CBA8",
		x"CBC3CBC2CBC1CBC0FFFFFFFFFFFFFFFFCBBFCBBECBBDCBBCCBBBCBBACBB9CBB8",
		x"CBD3CBD2CBD1CBD0CBCFCBCECBCDCBCCCBCBCBCACBC9CBC8CBC7CBC6CBC5CBC4",
		x"CBE3CBE2CBE1CBE0CBDFCBDECBDDCBDCCBDBCBDACBD9CBD8CBD7CBD6CBD5CBD4",
		x"CBF3CBF2CBF1CBF0CBEFCBEECBEDCBECCBEBCBEACBE9CBE8CBE7CBE6CBE5CBE4",
		x"FFFFFFFFFFFFFFFFCBFFCBFECBFDCBFCCBFBCBFACBF9CBF8CBF7CBF6CBF5CBF4",
		x"CC0FCC0ECC0DCC0CCC0BCC0ACC09CC08CC07CC06CC05CC04CC03CC02CC01CC00",
		x"CC1FCC1ECC1DCC1CCC1BCC1ACC19CC18CC17CC16CC15CC14CC13CC12CC11CC10",
		x"CC2FCC2ECC2DCC2CCC2BCC2ACC29CC28CC27CC26CC25CC24CC23CC22CC21CC20",
		x"CC3FCC3ECC3DCC3CCC3BCC3ACC39CC38CC37CC36CC35CC34CC33CC32CC31CC30",
		x"CC4BCC4ACC49CC48CC47CC46CC45CC44CC43CC42CC41CC40FFFFFFFFFFFFFFFF",
		x"CC5BCC5ACC59CC58CC57CC56CC55CC54CC53CC52CC51CC50CC4FCC4ECC4DCC4C",
		x"CC6BCC6ACC69CC68CC67CC66CC65CC64CC63CC62CC61CC60CC5FCC5ECC5DCC5C",
		x"CC7BCC7ACC79CC78CC77CC76CC75CC74CC73CC72CC71CC70CC6FCC6ECC6DCC6C",
		x"CC87CC86CC85CC84CC83CC82CC81CC80FFFFFFFFFFFFFFFFCC7FCC7ECC7DCC7C",
		x"CC97CC96CC95CC94CC93CC92CC91CC90CC8FCC8ECC8DCC8CCC8BCC8ACC89CC88",
		x"CCA7CCA6CCA5CCA4CCA3CCA2CCA1CCA0CC9FCC9ECC9DCC9CCC9BCC9ACC99CC98",
		x"CCB7CCB6CCB5CCB4CCB3CCB2CCB1CCB0CCAFCCAECCADCCACCCABCCAACCA9CCA8",
		x"CCC3CCC2CCC1CCC0FFFFFFFFFFFFFFFFCCBFCCBECCBDCCBCCCBBCCBACCB9CCB8",
		x"CCD3CCD2CCD1CCD0CCCFCCCECCCDCCCCCCCBCCCACCC9CCC8CCC7CCC6CCC5CCC4",
		x"CCE3CCE2CCE1CCE0CCDFCCDECCDDCCDCCCDBCCDACCD9CCD8CCD7CCD6CCD5CCD4",
		x"CCF3CCF2CCF1CCF0CCEFCCEECCEDCCECCCEBCCEACCE9CCE8CCE7CCE6CCE5CCE4",
		x"FFFFFFFFFFFFFFFFCCFFCCFECCFDCCFCCCFBCCFACCF9CCF8CCF7CCF6CCF5CCF4",
		x"CD0FCD0ECD0DCD0CCD0BCD0ACD09CD08CD07CD06CD05CD04CD03CD02CD01CD00",
		x"CD1FCD1ECD1DCD1CCD1BCD1ACD19CD18CD17CD16CD15CD14CD13CD12CD11CD10",
		x"CD2FCD2ECD2DCD2CCD2BCD2ACD29CD28CD27CD26CD25CD24CD23CD22CD21CD20",
		x"CD3FCD3ECD3DCD3CCD3BCD3ACD39CD38CD37CD36CD35CD34CD33CD32CD31CD30",
		x"CD4BCD4ACD49CD48CD47CD46CD45CD44CD43CD42CD41CD40FFFFFFFFFFFFFFFF",
		x"CD5BCD5ACD59CD58CD57CD56CD55CD54CD53CD52CD51CD50CD4FCD4ECD4DCD4C",
		x"CD6BCD6ACD69CD68CD67CD66CD65CD64CD63CD62CD61CD60CD5FCD5ECD5DCD5C",
		x"CD7BCD7ACD79CD78CD77CD76CD75CD74CD73CD72CD71CD70CD6FCD6ECD6DCD6C",
		x"CD87CD86CD85CD84CD83CD82CD81CD80FFFFFFFFFFFFFFFFCD7FCD7ECD7DCD7C",
		x"CD97CD96CD95CD94CD93CD92CD91CD90CD8FCD8ECD8DCD8CCD8BCD8ACD89CD88",
		x"CDA7CDA6CDA5CDA4CDA3CDA2CDA1CDA0CD9FCD9ECD9DCD9CCD9BCD9ACD99CD98",
		x"CDB7CDB6CDB5CDB4CDB3CDB2CDB1CDB0CDAFCDAECDADCDACCDABCDAACDA9CDA8",
		x"CDC3CDC2CDC1CDC0FFFFFFFFFFFFFFFFCDBFCDBECDBDCDBCCDBBCDBACDB9CDB8",
		x"CDD3CDD2CDD1CDD0CDCFCDCECDCDCDCCCDCBCDCACDC9CDC8CDC7CDC6CDC5CDC4",
		x"CDE3CDE2CDE1CDE0CDDFCDDECDDDCDDCCDDBCDDACDD9CDD8CDD7CDD6CDD5CDD4",
		x"CDF3CDF2CDF1CDF0CDEFCDEECDEDCDECCDEBCDEACDE9CDE8CDE7CDE6CDE5CDE4",
		x"FFFFFFFFFFFFFFFFCDFFCDFECDFDCDFCCDFBCDFACDF9CDF8CDF7CDF6CDF5CDF4",
		x"CE0FCE0ECE0DCE0CCE0BCE0ACE09CE08CE07CE06CE05CE04CE03CE02CE01CE00",
		x"CE1FCE1ECE1DCE1CCE1BCE1ACE19CE18CE17CE16CE15CE14CE13CE12CE11CE10",
		x"CE2FCE2ECE2DCE2CCE2BCE2ACE29CE28CE27CE26CE25CE24CE23CE22CE21CE20",
		x"CE3FCE3ECE3DCE3CCE3BCE3ACE39CE38CE37CE36CE35CE34CE33CE32CE31CE30",
		x"CE4BCE4ACE49CE48CE47CE46CE45CE44CE43CE42CE41CE40FFFFFFFFFFFFFFFF",
		x"CE5BCE5ACE59CE58CE57CE56CE55CE54CE53CE52CE51CE50CE4FCE4ECE4DCE4C",
		x"CE6BCE6ACE69CE68CE67CE66CE65CE64CE63CE62CE61CE60CE5FCE5ECE5DCE5C",
		x"CE7BCE7ACE79CE78CE77CE76CE75CE74CE73CE72CE71CE70CE6FCE6ECE6DCE6C",
		x"CE87CE86CE85CE84CE83CE82CE81CE80FFFFFFFFFFFFFFFFCE7FCE7ECE7DCE7C",
		x"CE97CE96CE95CE94CE93CE92CE91CE90CE8FCE8ECE8DCE8CCE8BCE8ACE89CE88",
		x"CEA7CEA6CEA5CEA4CEA3CEA2CEA1CEA0CE9FCE9ECE9DCE9CCE9BCE9ACE99CE98",
		x"CEB7CEB6CEB5CEB4CEB3CEB2CEB1CEB0CEAFCEAECEADCEACCEABCEAACEA9CEA8",
		x"CEC3CEC2CEC1CEC0FFFFFFFFFFFFFFFFCEBFCEBECEBDCEBCCEBBCEBACEB9CEB8",
		x"CED3CED2CED1CED0CECFCECECECDCECCCECBCECACEC9CEC8CEC7CEC6CEC5CEC4",
		x"CEE3CEE2CEE1CEE0CEDFCEDECEDDCEDCCEDBCEDACED9CED8CED7CED6CED5CED4",
		x"CEF3CEF2CEF1CEF0CEEFCEEECEEDCEECCEEBCEEACEE9CEE8CEE7CEE6CEE5CEE4",
		x"FFFFFFFFFFFFFFFFCEFFCEFECEFDCEFCCEFBCEFACEF9CEF8CEF7CEF6CEF5CEF4",
		x"CF0FCF0ECF0DCF0CCF0BCF0ACF09CF08CF07CF06CF05CF04CF03CF02CF01CF00",
		x"CF1FCF1ECF1DCF1CCF1BCF1ACF19CF18CF17CF16CF15CF14CF13CF12CF11CF10",
		x"CF2FCF2ECF2DCF2CCF2BCF2ACF29CF28CF27CF26CF25CF24CF23CF22CF21CF20",
		x"CF3FCF3ECF3DCF3CCF3BCF3ACF39CF38CF37CF36CF35CF34CF33CF32CF31CF30",
		x"CF4BCF4ACF49CF48CF47CF46CF45CF44CF43CF42CF41CF40FFFFFFFFFFFFFFFF",
		x"CF5BCF5ACF59CF58CF57CF56CF55CF54CF53CF52CF51CF50CF4FCF4ECF4DCF4C",
		x"CF6BCF6ACF69CF68CF67CF66CF65CF64CF63CF62CF61CF60CF5FCF5ECF5DCF5C",
		x"CF7BCF7ACF79CF78CF77CF76CF75CF74CF73CF72CF71CF70CF6FCF6ECF6DCF6C",
		x"CF87CF86CF85CF84CF83CF82CF81CF80FFFFFFFFFFFFFFFFCF7FCF7ECF7DCF7C",
		x"CF97CF96CF95CF94CF93CF92CF91CF90CF8FCF8ECF8DCF8CCF8BCF8ACF89CF88",
		x"CFA7CFA6CFA5CFA4CFA3CFA2CFA1CFA0CF9FCF9ECF9DCF9CCF9BCF9ACF99CF98",
		x"CFB7CFB6CFB5CFB4CFB3CFB2CFB1CFB0CFAFCFAECFADCFACCFABCFAACFA9CFA8",
		x"CFC3CFC2CFC1CFC0FFFFFFFFFFFFFFFFCFBFCFBECFBDCFBCCFBBCFBACFB9CFB8",
		x"CFD3CFD2CFD1CFD0CFCFCFCECFCDCFCCCFCBCFCACFC9CFC8CFC7CFC6CFC5CFC4",
		x"CFE3CFE2CFE1CFE0CFDFCFDECFDDCFDCCFDBCFDACFD9CFD8CFD7CFD6CFD5CFD4",
		x"CFF3CFF2CFF1CFF0CFEFCFEECFEDCFECCFEBCFEACFE9CFE8CFE7CFE6CFE5CFE4",
		x"FFFFFFFFFFFFFFFFCFFFCFFECFFDCFFCCFFBCFFACFF9CFF8CFF7CFF6CFF5CFF4",
		x"D00FD00ED00DD00CD00BD00AD009D008D007D006D005D004D003D002D001D000",
		x"D01FD01ED01DD01CD01BD01AD019D018D017D016D015D014D013D012D011D010",
		x"D02FD02ED02DD02CD02BD02AD029D028D027D026D025D024D023D022D021D020",
		x"D03FD03ED03DD03CD03BD03AD039D038D037D036D035D034D033D032D031D030",
		x"D04BD04AD049D048D047D046D045D044D043D042D041D040FFFFFFFFFFFFFFFF",
		x"D05BD05AD059D058D057D056D055D054D053D052D051D050D04FD04ED04DD04C",
		x"D06BD06AD069D068D067D066D065D064D063D062D061D060D05FD05ED05DD05C",
		x"D07BD07AD079D078D077D076D075D074D073D072D071D070D06FD06ED06DD06C",
		x"D087D086D085D084D083D082D081D080FFFFFFFFFFFFFFFFD07FD07ED07DD07C",
		x"D097D096D095D094D093D092D091D090D08FD08ED08DD08CD08BD08AD089D088",
		x"D0A7D0A6D0A5D0A4D0A3D0A2D0A1D0A0D09FD09ED09DD09CD09BD09AD099D098",
		x"D0B7D0B6D0B5D0B4D0B3D0B2D0B1D0B0D0AFD0AED0ADD0ACD0ABD0AAD0A9D0A8",
		x"D0C3D0C2D0C1D0C0FFFFFFFFFFFFFFFFD0BFD0BED0BDD0BCD0BBD0BAD0B9D0B8",
		x"D0D3D0D2D0D1D0D0D0CFD0CED0CDD0CCD0CBD0CAD0C9D0C8D0C7D0C6D0C5D0C4",
		x"D0E3D0E2D0E1D0E0D0DFD0DED0DDD0DCD0DBD0DAD0D9D0D8D0D7D0D6D0D5D0D4",
		x"D0F3D0F2D0F1D0F0D0EFD0EED0EDD0ECD0EBD0EAD0E9D0E8D0E7D0E6D0E5D0E4",
		x"FFFFFFFFFFFFFFFFD0FFD0FED0FDD0FCD0FBD0FAD0F9D0F8D0F7D0F6D0F5D0F4",
		x"D10FD10ED10DD10CD10BD10AD109D108D107D106D105D104D103D102D101D100",
		x"D11FD11ED11DD11CD11BD11AD119D118D117D116D115D114D113D112D111D110",
		x"D12FD12ED12DD12CD12BD12AD129D128D127D126D125D124D123D122D121D120",
		x"D13FD13ED13DD13CD13BD13AD139D138D137D136D135D134D133D132D131D130",
		x"D14BD14AD149D148D147D146D145D144D143D142D141D140FFFFFFFFFFFFFFFF",
		x"D15BD15AD159D158D157D156D155D154D153D152D151D150D14FD14ED14DD14C",
		x"D16BD16AD169D168D167D166D165D164D163D162D161D160D15FD15ED15DD15C",
		x"D17BD17AD179D178D177D176D175D174D173D172D171D170D16FD16ED16DD16C",
		x"D187D186D185D184D183D182D181D180FFFFFFFFFFFFFFFFD17FD17ED17DD17C",
		x"D197D196D195D194D193D192D191D190D18FD18ED18DD18CD18BD18AD189D188",
		x"D1A7D1A6D1A5D1A4D1A3D1A2D1A1D1A0D19FD19ED19DD19CD19BD19AD199D198",
		x"D1B7D1B6D1B5D1B4D1B3D1B2D1B1D1B0D1AFD1AED1ADD1ACD1ABD1AAD1A9D1A8",
		x"D1C3D1C2D1C1D1C0FFFFFFFFFFFFFFFFD1BFD1BED1BDD1BCD1BBD1BAD1B9D1B8",
		x"D1D3D1D2D1D1D1D0D1CFD1CED1CDD1CCD1CBD1CAD1C9D1C8D1C7D1C6D1C5D1C4",
		x"D1E3D1E2D1E1D1E0D1DFD1DED1DDD1DCD1DBD1DAD1D9D1D8D1D7D1D6D1D5D1D4",
		x"D1F3D1F2D1F1D1F0D1EFD1EED1EDD1ECD1EBD1EAD1E9D1E8D1E7D1E6D1E5D1E4",
		x"FFFFFFFFFFFFFFFFD1FFD1FED1FDD1FCD1FBD1FAD1F9D1F8D1F7D1F6D1F5D1F4",
		x"D20FD20ED20DD20CD20BD20AD209D208D207D206D205D204D203D202D201D200",
		x"D21FD21ED21DD21CD21BD21AD219D218D217D216D215D214D213D212D211D210",
		x"D22FD22ED22DD22CD22BD22AD229D228D227D226D225D224D223D222D221D220",
		x"D23FD23ED23DD23CD23BD23AD239D238D237D236D235D234D233D232D231D230",
		x"D24BD24AD249D248D247D246D245D244D243D242D241D240FFFFFFFFFFFFFFFF",
		x"D25BD25AD259D258D257D256D255D254D253D252D251D250D24FD24ED24DD24C",
		x"D26BD26AD269D268D267D266D265D264D263D262D261D260D25FD25ED25DD25C",
		x"D27BD27AD279D278D277D276D275D274D273D272D271D270D26FD26ED26DD26C",
		x"D287D286D285D284D283D282D281D280FFFFFFFFFFFFFFFFD27FD27ED27DD27C",
		x"D297D296D295D294D293D292D291D290D28FD28ED28DD28CD28BD28AD289D288",
		x"D2A7D2A6D2A5D2A4D2A3D2A2D2A1D2A0D29FD29ED29DD29CD29BD29AD299D298",
		x"D2B7D2B6D2B5D2B4D2B3D2B2D2B1D2B0D2AFD2AED2ADD2ACD2ABD2AAD2A9D2A8",
		x"D2C3D2C2D2C1D2C0FFFFFFFFFFFFFFFFD2BFD2BED2BDD2BCD2BBD2BAD2B9D2B8",
		x"D2D3D2D2D2D1D2D0D2CFD2CED2CDD2CCD2CBD2CAD2C9D2C8D2C7D2C6D2C5D2C4",
		x"D2E3D2E2D2E1D2E0D2DFD2DED2DDD2DCD2DBD2DAD2D9D2D8D2D7D2D6D2D5D2D4",
		x"D2F3D2F2D2F1D2F0D2EFD2EED2EDD2ECD2EBD2EAD2E9D2E8D2E7D2E6D2E5D2E4",
		x"FFFFFFFFFFFFFFFFD2FFD2FED2FDD2FCD2FBD2FAD2F9D2F8D2F7D2F6D2F5D2F4",
		x"D30FD30ED30DD30CD30BD30AD309D308D307D306D305D304D303D302D301D300",
		x"D31FD31ED31DD31CD31BD31AD319D318D317D316D315D314D313D312D311D310",
		x"D32FD32ED32DD32CD32BD32AD329D328D327D326D325D324D323D322D321D320",
		x"D33FD33ED33DD33CD33BD33AD339D338D337D336D335D334D333D332D331D330",
		x"D34BD34AD349D348D347D346D345D344D343D342D341D340FFFFFFFFFFFFFFFF",
		x"D35BD35AD359D358D357D356D355D354D353D352D351D350D34FD34ED34DD34C",
		x"D36BD36AD369D368D367D366D365D364D363D362D361D360D35FD35ED35DD35C",
		x"D37BD37AD379D378D377D376D375D374D373D372D371D370D36FD36ED36DD36C",
		x"D387D386D385D384D383D382D381D380FFFFFFFFFFFFFFFFD37FD37ED37DD37C",
		x"D397D396D395D394D393D392D391D390D38FD38ED38DD38CD38BD38AD389D388",
		x"D3A7D3A6D3A5D3A4D3A3D3A2D3A1D3A0D39FD39ED39DD39CD39BD39AD399D398",
		x"D3B7D3B6D3B5D3B4D3B3D3B2D3B1D3B0D3AFD3AED3ADD3ACD3ABD3AAD3A9D3A8",
		x"D3C3D3C2D3C1D3C0FFFFFFFFFFFFFFFFD3BFD3BED3BDD3BCD3BBD3BAD3B9D3B8",
		x"D3D3D3D2D3D1D3D0D3CFD3CED3CDD3CCD3CBD3CAD3C9D3C8D3C7D3C6D3C5D3C4",
		x"D3E3D3E2D3E1D3E0D3DFD3DED3DDD3DCD3DBD3DAD3D9D3D8D3D7D3D6D3D5D3D4",
		x"D3F3D3F2D3F1D3F0D3EFD3EED3EDD3ECD3EBD3EAD3E9D3E8D3E7D3E6D3E5D3E4",
		x"FFFFFFFFFFFFFFFFD3FFD3FED3FDD3FCD3FBD3FAD3F9D3F8D3F7D3F6D3F5D3F4",
		x"D40FD40ED40DD40CD40BD40AD409D408D407D406D405D404D403D402D401D400",
		x"D41FD41ED41DD41CD41BD41AD419D418D417D416D415D414D413D412D411D410",
		x"D42FD42ED42DD42CD42BD42AD429D428D427D426D425D424D423D422D421D420",
		x"D43FD43ED43DD43CD43BD43AD439D438D437D436D435D434D433D432D431D430",
		x"D44BD44AD449D448D447D446D445D444D443D442D441D440FFFFFFFFFFFFFFFF",
		x"D45BD45AD459D458D457D456D455D454D453D452D451D450D44FD44ED44DD44C",
		x"D46BD46AD469D468D467D466D465D464D463D462D461D460D45FD45ED45DD45C",
		x"D47BD47AD479D478D477D476D475D474D473D472D471D470D46FD46ED46DD46C",
		x"D487D486D485D484D483D482D481D480FFFFFFFFFFFFFFFFD47FD47ED47DD47C",
		x"D497D496D495D494D493D492D491D490D48FD48ED48DD48CD48BD48AD489D488",
		x"D4A7D4A6D4A5D4A4D4A3D4A2D4A1D4A0D49FD49ED49DD49CD49BD49AD499D498",
		x"D4B7D4B6D4B5D4B4D4B3D4B2D4B1D4B0D4AFD4AED4ADD4ACD4ABD4AAD4A9D4A8",
		x"D4C3D4C2D4C1D4C0FFFFFFFFFFFFFFFFD4BFD4BED4BDD4BCD4BBD4BAD4B9D4B8",
		x"D4D3D4D2D4D1D4D0D4CFD4CED4CDD4CCD4CBD4CAD4C9D4C8D4C7D4C6D4C5D4C4",
		x"D4E3D4E2D4E1D4E0D4DFD4DED4DDD4DCD4DBD4DAD4D9D4D8D4D7D4D6D4D5D4D4",
		x"D4F3D4F2D4F1D4F0D4EFD4EED4EDD4ECD4EBD4EAD4E9D4E8D4E7D4E6D4E5D4E4",
		x"FFFFFFFFFFFFFFFFD4FFD4FED4FDD4FCD4FBD4FAD4F9D4F8D4F7D4F6D4F5D4F4",
		x"D50FD50ED50DD50CD50BD50AD509D508D507D506D505D504D503D502D501D500",
		x"D51FD51ED51DD51CD51BD51AD519D518D517D516D515D514D513D512D511D510",
		x"D52FD52ED52DD52CD52BD52AD529D528D527D526D525D524D523D522D521D520",
		x"D53FD53ED53DD53CD53BD53AD539D538D537D536D535D534D533D532D531D530",
		x"D54BD54AD549D548D547D546D545D544D543D542D541D540FFFFFFFFFFFFFFFF",
		x"D55BD55AD559D558D557D556D555D554D553D552D551D550D54FD54ED54DD54C",
		x"D56BD56AD569D568D567D566D565D564D563D562D561D560D55FD55ED55DD55C",
		x"D57BD57AD579D578D577D576D575D574D573D572D571D570D56FD56ED56DD56C",
		x"D587D586D585D584D583D582D581D580FFFFFFFFFFFFFFFFD57FD57ED57DD57C",
		x"D597D596D595D594D593D592D591D590D58FD58ED58DD58CD58BD58AD589D588",
		x"D5A7D5A6D5A5D5A4D5A3D5A2D5A1D5A0D59FD59ED59DD59CD59BD59AD599D598",
		x"D5B7D5B6D5B5D5B4D5B3D5B2D5B1D5B0D5AFD5AED5ADD5ACD5ABD5AAD5A9D5A8",
		x"D5C3D5C2D5C1D5C0FFFFFFFFFFFFFFFFD5BFD5BED5BDD5BCD5BBD5BAD5B9D5B8",
		x"D5D3D5D2D5D1D5D0D5CFD5CED5CDD5CCD5CBD5CAD5C9D5C8D5C7D5C6D5C5D5C4",
		x"D5E3D5E2D5E1D5E0D5DFD5DED5DDD5DCD5DBD5DAD5D9D5D8D5D7D5D6D5D5D5D4",
		x"D5F3D5F2D5F1D5F0D5EFD5EED5EDD5ECD5EBD5EAD5E9D5E8D5E7D5E6D5E5D5E4",
		x"FFFFFFFFFFFFFFFFD5FFD5FED5FDD5FCD5FBD5FAD5F9D5F8D5F7D5F6D5F5D5F4",
		x"D60FD60ED60DD60CD60BD60AD609D608D607D606D605D604D603D602D601D600",
		x"D61FD61ED61DD61CD61BD61AD619D618D617D616D615D614D613D612D611D610",
		x"D62FD62ED62DD62CD62BD62AD629D628D627D626D625D624D623D622D621D620",
		x"D63FD63ED63DD63CD63BD63AD639D638D637D636D635D634D633D632D631D630",
		x"D64BD64AD649D648D647D646D645D644D643D642D641D640FFFFFFFFFFFFFFFF",
		x"D65BD65AD659D658D657D656D655D654D653D652D651D650D64FD64ED64DD64C",
		x"D66BD66AD669D668D667D666D665D664D663D662D661D660D65FD65ED65DD65C",
		x"D67BD67AD679D678D677D676D675D674D673D672D671D670D66FD66ED66DD66C",
		x"D687D686D685D684D683D682D681D680FFFFFFFFFFFFFFFFD67FD67ED67DD67C",
		x"D697D696D695D694D693D692D691D690D68FD68ED68DD68CD68BD68AD689D688",
		x"D6A7D6A6D6A5D6A4D6A3D6A2D6A1D6A0D69FD69ED69DD69CD69BD69AD699D698",
		x"D6B7D6B6D6B5D6B4D6B3D6B2D6B1D6B0D6AFD6AED6ADD6ACD6ABD6AAD6A9D6A8",
		x"D6C3D6C2D6C1D6C0FFFFFFFFFFFFFFFFD6BFD6BED6BDD6BCD6BBD6BAD6B9D6B8",
		x"D6D3D6D2D6D1D6D0D6CFD6CED6CDD6CCD6CBD6CAD6C9D6C8D6C7D6C6D6C5D6C4",
		x"D6E3D6E2D6E1D6E0D6DFD6DED6DDD6DCD6DBD6DAD6D9D6D8D6D7D6D6D6D5D6D4",
		x"D6F3D6F2D6F1D6F0D6EFD6EED6EDD6ECD6EBD6EAD6E9D6E8D6E7D6E6D6E5D6E4",
		x"FFFFFFFFFFFFFFFFD6FFD6FED6FDD6FCD6FBD6FAD6F9D6F8D6F7D6F6D6F5D6F4",
		x"D70FD70ED70DD70CD70BD70AD709D708D707D706D705D704D703D702D701D700",
		x"D71FD71ED71DD71CD71BD71AD719D718D717D716D715D714D713D712D711D710",
		x"D72FD72ED72DD72CD72BD72AD729D728D727D726D725D724D723D722D721D720",
		x"D73FD73ED73DD73CD73BD73AD739D738D737D736D735D734D733D732D731D730",
		x"D74BD74AD749D748D747D746D745D744D743D742D741D740FFFFFFFFFFFFFFFF",
		x"D75BD75AD759D758D757D756D755D754D753D752D751D750D74FD74ED74DD74C",
		x"D76BD76AD769D768D767D766D765D764D763D762D761D760D75FD75ED75DD75C",
		x"D77BD77AD779D778D777D776D775D774D773D772D771D770D76FD76ED76DD76C",
		x"D787D786D785D784D783D782D781D780FFFFFFFFFFFFFFFFD77FD77ED77DD77C",
		x"D797D796D795D794D793D792D791D790D78FD78ED78DD78CD78BD78AD789D788",
		x"D7A7D7A6D7A5D7A4D7A3D7A2D7A1D7A0D79FD79ED79DD79CD79BD79AD799D798",
		x"D7B7D7B6D7B5D7B4D7B3D7B2D7B1D7B0D7AFD7AED7ADD7ACD7ABD7AAD7A9D7A8",
		x"D7C3D7C2D7C1D7C0FFFFFFFFFFFFFFFFD7BFD7BED7BDD7BCD7BBD7BAD7B9D7B8",
		x"D7D3D7D2D7D1D7D0D7CFD7CED7CDD7CCD7CBD7CAD7C9D7C8D7C7D7C6D7C5D7C4",
		x"D7E3D7E2D7E1D7E0D7DFD7DED7DDD7DCD7DBD7DAD7D9D7D8D7D7D7D6D7D5D7D4",
		x"D7F3D7F2D7F1D7F0D7EFD7EED7EDD7ECD7EBD7EAD7E9D7E8D7E7D7E6D7E5D7E4",
		x"FFFFFFFFFFFFFFFFD7FFD7FED7FDD7FCD7FBD7FAD7F9D7F8D7F7D7F6D7F5D7F4",
		x"D80FD80ED80DD80CD80BD80AD809D808D807D806D805D804D803D802D801D800",
		x"D81FD81ED81DD81CD81BD81AD819D818D817D816D815D814D813D812D811D810",
		x"D82FD82ED82DD82CD82BD82AD829D828D827D826D825D824D823D822D821D820",
		x"D83FD83ED83DD83CD83BD83AD839D838D837D836D835D834D833D832D831D830",
		x"D84BD84AD849D848D847D846D845D844D843D842D841D840FFFFFFFFFFFFFFFF",
		x"D85BD85AD859D858D857D856D855D854D853D852D851D850D84FD84ED84DD84C",
		x"D86BD86AD869D868D867D866D865D864D863D862D861D860D85FD85ED85DD85C",
		x"D87BD87AD879D878D877D876D875D874D873D872D871D870D86FD86ED86DD86C",
		x"D887D886D885D884D883D882D881D880FFFFFFFFFFFFFFFFD87FD87ED87DD87C",
		x"D897D896D895D894D893D892D891D890D88FD88ED88DD88CD88BD88AD889D888",
		x"D8A7D8A6D8A5D8A4D8A3D8A2D8A1D8A0D89FD89ED89DD89CD89BD89AD899D898",
		x"D8B7D8B6D8B5D8B4D8B3D8B2D8B1D8B0D8AFD8AED8ADD8ACD8ABD8AAD8A9D8A8",
		x"D8C3D8C2D8C1D8C0FFFFFFFFFFFFFFFFD8BFD8BED8BDD8BCD8BBD8BAD8B9D8B8",
		x"D8D3D8D2D8D1D8D0D8CFD8CED8CDD8CCD8CBD8CAD8C9D8C8D8C7D8C6D8C5D8C4",
		x"D8E3D8E2D8E1D8E0D8DFD8DED8DDD8DCD8DBD8DAD8D9D8D8D8D7D8D6D8D5D8D4",
		x"D8F3D8F2D8F1D8F0D8EFD8EED8EDD8ECD8EBD8EAD8E9D8E8D8E7D8E6D8E5D8E4",
		x"FFFFFFFFFFFFFFFFD8FFD8FED8FDD8FCD8FBD8FAD8F9D8F8D8F7D8F6D8F5D8F4",
		x"D90FD90ED90DD90CD90BD90AD909D908D907D906D905D904D903D902D901D900",
		x"D91FD91ED91DD91CD91BD91AD919D918D917D916D915D914D913D912D911D910",
		x"D92FD92ED92DD92CD92BD92AD929D928D927D926D925D924D923D922D921D920",
		x"D93FD93ED93DD93CD93BD93AD939D938D937D936D935D934D933D932D931D930",
		x"D94BD94AD949D948D947D946D945D944D943D942D941D940FFFFFFFFFFFFFFFF",
		x"D95BD95AD959D958D957D956D955D954D953D952D951D950D94FD94ED94DD94C",
		x"D96BD96AD969D968D967D966D965D964D963D962D961D960D95FD95ED95DD95C",
		x"D97BD97AD979D978D977D976D975D974D973D972D971D970D96FD96ED96DD96C",
		x"D987D986D985D984D983D982D981D980FFFFFFFFFFFFFFFFD97FD97ED97DD97C",
		x"D997D996D995D994D993D992D991D990D98FD98ED98DD98CD98BD98AD989D988",
		x"D9A7D9A6D9A5D9A4D9A3D9A2D9A1D9A0D99FD99ED99DD99CD99BD99AD999D998",
		x"D9B7D9B6D9B5D9B4D9B3D9B2D9B1D9B0D9AFD9AED9ADD9ACD9ABD9AAD9A9D9A8",
		x"D9C3D9C2D9C1D9C0FFFFFFFFFFFFFFFFD9BFD9BED9BDD9BCD9BBD9BAD9B9D9B8",
		x"D9D3D9D2D9D1D9D0D9CFD9CED9CDD9CCD9CBD9CAD9C9D9C8D9C7D9C6D9C5D9C4",
		x"D9E3D9E2D9E1D9E0D9DFD9DED9DDD9DCD9DBD9DAD9D9D9D8D9D7D9D6D9D5D9D4",
		x"D9F3D9F2D9F1D9F0D9EFD9EED9EDD9ECD9EBD9EAD9E9D9E8D9E7D9E6D9E5D9E4",
		x"FFFFFFFFFFFFFFFFD9FFD9FED9FDD9FCD9FBD9FAD9F9D9F8D9F7D9F6D9F5D9F4",
		x"DA0FDA0EDA0DDA0CDA0BDA0ADA09DA08DA07DA06DA05DA04DA03DA02DA01DA00",
		x"DA1FDA1EDA1DDA1CDA1BDA1ADA19DA18DA17DA16DA15DA14DA13DA12DA11DA10",
		x"DA2FDA2EDA2DDA2CDA2BDA2ADA29DA28DA27DA26DA25DA24DA23DA22DA21DA20",
		x"DA3FDA3EDA3DDA3CDA3BDA3ADA39DA38DA37DA36DA35DA34DA33DA32DA31DA30",
		x"DA4BDA4ADA49DA48DA47DA46DA45DA44DA43DA42DA41DA40FFFFFFFFFFFFFFFF",
		x"DA5BDA5ADA59DA58DA57DA56DA55DA54DA53DA52DA51DA50DA4FDA4EDA4DDA4C",
		x"DA6BDA6ADA69DA68DA67DA66DA65DA64DA63DA62DA61DA60DA5FDA5EDA5DDA5C",
		x"DA7BDA7ADA79DA78DA77DA76DA75DA74DA73DA72DA71DA70DA6FDA6EDA6DDA6C",
		x"DA87DA86DA85DA84DA83DA82DA81DA80FFFFFFFFFFFFFFFFDA7FDA7EDA7DDA7C",
		x"DA97DA96DA95DA94DA93DA92DA91DA90DA8FDA8EDA8DDA8CDA8BDA8ADA89DA88",
		x"DAA7DAA6DAA5DAA4DAA3DAA2DAA1DAA0DA9FDA9EDA9DDA9CDA9BDA9ADA99DA98",
		x"DAB7DAB6DAB5DAB4DAB3DAB2DAB1DAB0DAAFDAAEDAADDAACDAABDAAADAA9DAA8",
		x"DAC3DAC2DAC1DAC0FFFFFFFFFFFFFFFFDABFDABEDABDDABCDABBDABADAB9DAB8",
		x"DAD3DAD2DAD1DAD0DACFDACEDACDDACCDACBDACADAC9DAC8DAC7DAC6DAC5DAC4",
		x"DAE3DAE2DAE1DAE0DADFDADEDADDDADCDADBDADADAD9DAD8DAD7DAD6DAD5DAD4",
		x"DAF3DAF2DAF1DAF0DAEFDAEEDAEDDAECDAEBDAEADAE9DAE8DAE7DAE6DAE5DAE4",
		x"FFFFFFFFFFFFFFFFDAFFDAFEDAFDDAFCDAFBDAFADAF9DAF8DAF7DAF6DAF5DAF4",
		x"DB0FDB0EDB0DDB0CDB0BDB0ADB09DB08DB07DB06DB05DB04DB03DB02DB01DB00",
		x"DB1FDB1EDB1DDB1CDB1BDB1ADB19DB18DB17DB16DB15DB14DB13DB12DB11DB10",
		x"DB2FDB2EDB2DDB2CDB2BDB2ADB29DB28DB27DB26DB25DB24DB23DB22DB21DB20",
		x"DB3FDB3EDB3DDB3CDB3BDB3ADB39DB38DB37DB36DB35DB34DB33DB32DB31DB30",
		x"DB4BDB4ADB49DB48DB47DB46DB45DB44DB43DB42DB41DB40FFFFFFFFFFFFFFFF",
		x"DB5BDB5ADB59DB58DB57DB56DB55DB54DB53DB52DB51DB50DB4FDB4EDB4DDB4C",
		x"DB6BDB6ADB69DB68DB67DB66DB65DB64DB63DB62DB61DB60DB5FDB5EDB5DDB5C",
		x"DB7BDB7ADB79DB78DB77DB76DB75DB74DB73DB72DB71DB70DB6FDB6EDB6DDB6C",
		x"DB87DB86DB85DB84DB83DB82DB81DB80FFFFFFFFFFFFFFFFDB7FDB7EDB7DDB7C",
		x"DB97DB96DB95DB94DB93DB92DB91DB90DB8FDB8EDB8DDB8CDB8BDB8ADB89DB88",
		x"DBA7DBA6DBA5DBA4DBA3DBA2DBA1DBA0DB9FDB9EDB9DDB9CDB9BDB9ADB99DB98",
		x"DBB7DBB6DBB5DBB4DBB3DBB2DBB1DBB0DBAFDBAEDBADDBACDBABDBAADBA9DBA8",
		x"DBC3DBC2DBC1DBC0FFFFFFFFFFFFFFFFDBBFDBBEDBBDDBBCDBBBDBBADBB9DBB8",
		x"DBD3DBD2DBD1DBD0DBCFDBCEDBCDDBCCDBCBDBCADBC9DBC8DBC7DBC6DBC5DBC4",
		x"DBE3DBE2DBE1DBE0DBDFDBDEDBDDDBDCDBDBDBDADBD9DBD8DBD7DBD6DBD5DBD4",
		x"DBF3DBF2DBF1DBF0DBEFDBEEDBEDDBECDBEBDBEADBE9DBE8DBE7DBE6DBE5DBE4",
		x"FFFFFFFFFFFFFFFFDBFFDBFEDBFDDBFCDBFBDBFADBF9DBF8DBF7DBF6DBF5DBF4",
		x"DC0FDC0EDC0DDC0CDC0BDC0ADC09DC08DC07DC06DC05DC04DC03DC02DC01DC00",
		x"DC1FDC1EDC1DDC1CDC1BDC1ADC19DC18DC17DC16DC15DC14DC13DC12DC11DC10",
		x"DC2FDC2EDC2DDC2CDC2BDC2ADC29DC28DC27DC26DC25DC24DC23DC22DC21DC20",
		x"DC3FDC3EDC3DDC3CDC3BDC3ADC39DC38DC37DC36DC35DC34DC33DC32DC31DC30",
		x"DC4BDC4ADC49DC48DC47DC46DC45DC44DC43DC42DC41DC40FFFFFFFFFFFFFFFF",
		x"DC5BDC5ADC59DC58DC57DC56DC55DC54DC53DC52DC51DC50DC4FDC4EDC4DDC4C",
		x"DC6BDC6ADC69DC68DC67DC66DC65DC64DC63DC62DC61DC60DC5FDC5EDC5DDC5C",
		x"DC7BDC7ADC79DC78DC77DC76DC75DC74DC73DC72DC71DC70DC6FDC6EDC6DDC6C",
		x"DC87DC86DC85DC84DC83DC82DC81DC80FFFFFFFFFFFFFFFFDC7FDC7EDC7DDC7C",
		x"DC97DC96DC95DC94DC93DC92DC91DC90DC8FDC8EDC8DDC8CDC8BDC8ADC89DC88",
		x"DCA7DCA6DCA5DCA4DCA3DCA2DCA1DCA0DC9FDC9EDC9DDC9CDC9BDC9ADC99DC98",
		x"DCB7DCB6DCB5DCB4DCB3DCB2DCB1DCB0DCAFDCAEDCADDCACDCABDCAADCA9DCA8",
		x"DCC3DCC2DCC1DCC0FFFFFFFFFFFFFFFFDCBFDCBEDCBDDCBCDCBBDCBADCB9DCB8",
		x"DCD3DCD2DCD1DCD0DCCFDCCEDCCDDCCCDCCBDCCADCC9DCC8DCC7DCC6DCC5DCC4",
		x"DCE3DCE2DCE1DCE0DCDFDCDEDCDDDCDCDCDBDCDADCD9DCD8DCD7DCD6DCD5DCD4",
		x"DCF3DCF2DCF1DCF0DCEFDCEEDCEDDCECDCEBDCEADCE9DCE8DCE7DCE6DCE5DCE4",
		x"FFFFFFFFFFFFFFFFDCFFDCFEDCFDDCFCDCFBDCFADCF9DCF8DCF7DCF6DCF5DCF4",
		x"DD0FDD0EDD0DDD0CDD0BDD0ADD09DD08DD07DD06DD05DD04DD03DD02DD01DD00",
		x"DD1FDD1EDD1DDD1CDD1BDD1ADD19DD18DD17DD16DD15DD14DD13DD12DD11DD10",
		x"DD2FDD2EDD2DDD2CDD2BDD2ADD29DD28DD27DD26DD25DD24DD23DD22DD21DD20",
		x"DD3FDD3EDD3DDD3CDD3BDD3ADD39DD38DD37DD36DD35DD34DD33DD32DD31DD30",
		x"DD4BDD4ADD49DD48DD47DD46DD45DD44DD43DD42DD41DD40FFFFFFFFFFFFFFFF",
		x"DD5BDD5ADD59DD58DD57DD56DD55DD54DD53DD52DD51DD50DD4FDD4EDD4DDD4C",
		x"DD6BDD6ADD69DD68DD67DD66DD65DD64DD63DD62DD61DD60DD5FDD5EDD5DDD5C",
		x"DD7BDD7ADD79DD78DD77DD76DD75DD74DD73DD72DD71DD70DD6FDD6EDD6DDD6C",
		x"DD87DD86DD85DD84DD83DD82DD81DD80FFFFFFFFFFFFFFFFDD7FDD7EDD7DDD7C",
		x"DD97DD96DD95DD94DD93DD92DD91DD90DD8FDD8EDD8DDD8CDD8BDD8ADD89DD88",
		x"DDA7DDA6DDA5DDA4DDA3DDA2DDA1DDA0DD9FDD9EDD9DDD9CDD9BDD9ADD99DD98",
		x"DDB7DDB6DDB5DDB4DDB3DDB2DDB1DDB0DDAFDDAEDDADDDACDDABDDAADDA9DDA8",
		x"DDC3DDC2DDC1DDC0FFFFFFFFFFFFFFFFDDBFDDBEDDBDDDBCDDBBDDBADDB9DDB8",
		x"DDD3DDD2DDD1DDD0DDCFDDCEDDCDDDCCDDCBDDCADDC9DDC8DDC7DDC6DDC5DDC4",
		x"DDE3DDE2DDE1DDE0DDDFDDDEDDDDDDDCDDDBDDDADDD9DDD8DDD7DDD6DDD5DDD4",
		x"DDF3DDF2DDF1DDF0DDEFDDEEDDEDDDECDDEBDDEADDE9DDE8DDE7DDE6DDE5DDE4",
		x"FFFFFFFFFFFFFFFFDDFFDDFEDDFDDDFCDDFBDDFADDF9DDF8DDF7DDF6DDF5DDF4",
		x"DE0FDE0EDE0DDE0CDE0BDE0ADE09DE08DE07DE06DE05DE04DE03DE02DE01DE00",
		x"DE1FDE1EDE1DDE1CDE1BDE1ADE19DE18DE17DE16DE15DE14DE13DE12DE11DE10",
		x"DE2FDE2EDE2DDE2CDE2BDE2ADE29DE28DE27DE26DE25DE24DE23DE22DE21DE20",
		x"DE3FDE3EDE3DDE3CDE3BDE3ADE39DE38DE37DE36DE35DE34DE33DE32DE31DE30",
		x"DE4BDE4ADE49DE48DE47DE46DE45DE44DE43DE42DE41DE40FFFFFFFFFFFFFFFF",
		x"DE5BDE5ADE59DE58DE57DE56DE55DE54DE53DE52DE51DE50DE4FDE4EDE4DDE4C",
		x"DE6BDE6ADE69DE68DE67DE66DE65DE64DE63DE62DE61DE60DE5FDE5EDE5DDE5C",
		x"DE7BDE7ADE79DE78DE77DE76DE75DE74DE73DE72DE71DE70DE6FDE6EDE6DDE6C",
		x"DE87DE86DE85DE84DE83DE82DE81DE80FFFFFFFFFFFFFFFFDE7FDE7EDE7DDE7C",
		x"DE97DE96DE95DE94DE93DE92DE91DE90DE8FDE8EDE8DDE8CDE8BDE8ADE89DE88",
		x"DEA7DEA6DEA5DEA4DEA3DEA2DEA1DEA0DE9FDE9EDE9DDE9CDE9BDE9ADE99DE98",
		x"DEB7DEB6DEB5DEB4DEB3DEB2DEB1DEB0DEAFDEAEDEADDEACDEABDEAADEA9DEA8",
		x"DEC3DEC2DEC1DEC0FFFFFFFFFFFFFFFFDEBFDEBEDEBDDEBCDEBBDEBADEB9DEB8",
		x"DED3DED2DED1DED0DECFDECEDECDDECCDECBDECADEC9DEC8DEC7DEC6DEC5DEC4",
		x"DEE3DEE2DEE1DEE0DEDFDEDEDEDDDEDCDEDBDEDADED9DED8DED7DED6DED5DED4",
		x"DEF3DEF2DEF1DEF0DEEFDEEEDEEDDEECDEEBDEEADEE9DEE8DEE7DEE6DEE5DEE4",
		x"FFFFFFFFFFFFFFFFDEFFDEFEDEFDDEFCDEFBDEFADEF9DEF8DEF7DEF6DEF5DEF4",
		x"DF0FDF0EDF0DDF0CDF0BDF0ADF09DF08DF07DF06DF05DF04DF03DF02DF01DF00",
		x"DF1FDF1EDF1DDF1CDF1BDF1ADF19DF18DF17DF16DF15DF14DF13DF12DF11DF10",
		x"DF2FDF2EDF2DDF2CDF2BDF2ADF29DF28DF27DF26DF25DF24DF23DF22DF21DF20",
		x"DF3FDF3EDF3DDF3CDF3BDF3ADF39DF38DF37DF36DF35DF34DF33DF32DF31DF30",
		x"DF4BDF4ADF49DF48DF47DF46DF45DF44DF43DF42DF41DF40FFFFFFFFFFFFFFFF",
		x"DF5BDF5ADF59DF58DF57DF56DF55DF54DF53DF52DF51DF50DF4FDF4EDF4DDF4C",
		x"DF6BDF6ADF69DF68DF67DF66DF65DF64DF63DF62DF61DF60DF5FDF5EDF5DDF5C",
		x"DF7BDF7ADF79DF78DF77DF76DF75DF74DF73DF72DF71DF70DF6FDF6EDF6DDF6C",
		x"DF87DF86DF85DF84DF83DF82DF81DF80FFFFFFFFFFFFFFFFDF7FDF7EDF7DDF7C",
		x"DF97DF96DF95DF94DF93DF92DF91DF90DF8FDF8EDF8DDF8CDF8BDF8ADF89DF88",
		x"DFA7DFA6DFA5DFA4DFA3DFA2DFA1DFA0DF9FDF9EDF9DDF9CDF9BDF9ADF99DF98",
		x"DFB7DFB6DFB5DFB4DFB3DFB2DFB1DFB0DFAFDFAEDFADDFACDFABDFAADFA9DFA8",
		x"DFC3DFC2DFC1DFC0FFFFFFFFFFFFFFFFDFBFDFBEDFBDDFBCDFBBDFBADFB9DFB8",
		x"DFD3DFD2DFD1DFD0DFCFDFCEDFCDDFCCDFCBDFCADFC9DFC8DFC7DFC6DFC5DFC4",
		x"DFE3DFE2DFE1DFE0DFDFDFDEDFDDDFDCDFDBDFDADFD9DFD8DFD7DFD6DFD5DFD4",
		x"DFF3DFF2DFF1DFF0DFEFDFEEDFEDDFECDFEBDFEADFE9DFE8DFE7DFE6DFE5DFE4",
		x"FFFFFFFFFFFFFFFFDFFFDFFEDFFDDFFCDFFBDFFADFF9DFF8DFF7DFF6DFF5DFF4",
		x"E00FE00EE00DE00CE00BE00AE009E008E007E006E005E004E003E002E001E000",
		x"E01FE01EE01DE01CE01BE01AE019E018E017E016E015E014E013E012E011E010",
		x"E02FE02EE02DE02CE02BE02AE029E028E027E026E025E024E023E022E021E020",
		x"E03FE03EE03DE03CE03BE03AE039E038E037E036E035E034E033E032E031E030",
		x"E04BE04AE049E048E047E046E045E044E043E042E041E040FFFFFFFFFFFFFFFF",
		x"E05BE05AE059E058E057E056E055E054E053E052E051E050E04FE04EE04DE04C",
		x"E06BE06AE069E068E067E066E065E064E063E062E061E060E05FE05EE05DE05C",
		x"E07BE07AE079E078E077E076E075E074E073E072E071E070E06FE06EE06DE06C",
		x"E087E086E085E084E083E082E081E080FFFFFFFFFFFFFFFFE07FE07EE07DE07C",
		x"E097E096E095E094E093E092E091E090E08FE08EE08DE08CE08BE08AE089E088",
		x"E0A7E0A6E0A5E0A4E0A3E0A2E0A1E0A0E09FE09EE09DE09CE09BE09AE099E098",
		x"E0B7E0B6E0B5E0B4E0B3E0B2E0B1E0B0E0AFE0AEE0ADE0ACE0ABE0AAE0A9E0A8",
		x"E0C3E0C2E0C1E0C0FFFFFFFFFFFFFFFFE0BFE0BEE0BDE0BCE0BBE0BAE0B9E0B8",
		x"E0D3E0D2E0D1E0D0E0CFE0CEE0CDE0CCE0CBE0CAE0C9E0C8E0C7E0C6E0C5E0C4",
		x"E0E3E0E2E0E1E0E0E0DFE0DEE0DDE0DCE0DBE0DAE0D9E0D8E0D7E0D6E0D5E0D4",
		x"E0F3E0F2E0F1E0F0E0EFE0EEE0EDE0ECE0EBE0EAE0E9E0E8E0E7E0E6E0E5E0E4",
		x"FFFFFFFFFFFFFFFFE0FFE0FEE0FDE0FCE0FBE0FAE0F9E0F8E0F7E0F6E0F5E0F4",
		x"E10FE10EE10DE10CE10BE10AE109E108E107E106E105E104E103E102E101E100",
		x"E11FE11EE11DE11CE11BE11AE119E118E117E116E115E114E113E112E111E110",
		x"E12FE12EE12DE12CE12BE12AE129E128E127E126E125E124E123E122E121E120",
		x"E13FE13EE13DE13CE13BE13AE139E138E137E136E135E134E133E132E131E130",
		x"E14BE14AE149E148E147E146E145E144E143E142E141E140FFFFFFFFFFFFFFFF",
		x"E15BE15AE159E158E157E156E155E154E153E152E151E150E14FE14EE14DE14C",
		x"E16BE16AE169E168E167E166E165E164E163E162E161E160E15FE15EE15DE15C",
		x"E17BE17AE179E178E177E176E175E174E173E172E171E170E16FE16EE16DE16C",
		x"E187E186E185E184E183E182E181E180FFFFFFFFFFFFFFFFE17FE17EE17DE17C",
		x"E197E196E195E194E193E192E191E190E18FE18EE18DE18CE18BE18AE189E188",
		x"E1A7E1A6E1A5E1A4E1A3E1A2E1A1E1A0E19FE19EE19DE19CE19BE19AE199E198",
		x"E1B7E1B6E1B5E1B4E1B3E1B2E1B1E1B0E1AFE1AEE1ADE1ACE1ABE1AAE1A9E1A8",
		x"E1C3E1C2E1C1E1C0FFFFFFFFFFFFFFFFE1BFE1BEE1BDE1BCE1BBE1BAE1B9E1B8",
		x"E1D3E1D2E1D1E1D0E1CFE1CEE1CDE1CCE1CBE1CAE1C9E1C8E1C7E1C6E1C5E1C4",
		x"E1E3E1E2E1E1E1E0E1DFE1DEE1DDE1DCE1DBE1DAE1D9E1D8E1D7E1D6E1D5E1D4",
		x"E1F3E1F2E1F1E1F0E1EFE1EEE1EDE1ECE1EBE1EAE1E9E1E8E1E7E1E6E1E5E1E4",
		x"FFFFFFFFFFFFFFFFE1FFE1FEE1FDE1FCE1FBE1FAE1F9E1F8E1F7E1F6E1F5E1F4",
		x"E20FE20EE20DE20CE20BE20AE209E208E207E206E205E204E203E202E201E200",
		x"E21FE21EE21DE21CE21BE21AE219E218E217E216E215E214E213E212E211E210",
		x"E22FE22EE22DE22CE22BE22AE229E228E227E226E225E224E223E222E221E220",
		x"E23FE23EE23DE23CE23BE23AE239E238E237E236E235E234E233E232E231E230",
		x"E24BE24AE249E248E247E246E245E244E243E242E241E240FFFFFFFFFFFFFFFF",
		x"E25BE25AE259E258E257E256E255E254E253E252E251E250E24FE24EE24DE24C",
		x"E26BE26AE269E268E267E266E265E264E263E262E261E260E25FE25EE25DE25C",
		x"E27BE27AE279E278E277E276E275E274E273E272E271E270E26FE26EE26DE26C",
		x"E287E286E285E284E283E282E281E280FFFFFFFFFFFFFFFFE27FE27EE27DE27C",
		x"E297E296E295E294E293E292E291E290E28FE28EE28DE28CE28BE28AE289E288",
		x"E2A7E2A6E2A5E2A4E2A3E2A2E2A1E2A0E29FE29EE29DE29CE29BE29AE299E298",
		x"E2B7E2B6E2B5E2B4E2B3E2B2E2B1E2B0E2AFE2AEE2ADE2ACE2ABE2AAE2A9E2A8",
		x"E2C3E2C2E2C1E2C0FFFFFFFFFFFFFFFFE2BFE2BEE2BDE2BCE2BBE2BAE2B9E2B8",
		x"E2D3E2D2E2D1E2D0E2CFE2CEE2CDE2CCE2CBE2CAE2C9E2C8E2C7E2C6E2C5E2C4",
		x"E2E3E2E2E2E1E2E0E2DFE2DEE2DDE2DCE2DBE2DAE2D9E2D8E2D7E2D6E2D5E2D4",
		x"E2F3E2F2E2F1E2F0E2EFE2EEE2EDE2ECE2EBE2EAE2E9E2E8E2E7E2E6E2E5E2E4",
		x"FFFFFFFFFFFFFFFFE2FFE2FEE2FDE2FCE2FBE2FAE2F9E2F8E2F7E2F6E2F5E2F4",
		x"E30FE30EE30DE30CE30BE30AE309E308E307E306E305E304E303E302E301E300",
		x"E31FE31EE31DE31CE31BE31AE319E318E317E316E315E314E313E312E311E310",
		x"E32FE32EE32DE32CE32BE32AE329E328E327E326E325E324E323E322E321E320",
		x"E33FE33EE33DE33CE33BE33AE339E338E337E336E335E334E333E332E331E330",
		x"E34BE34AE349E348E347E346E345E344E343E342E341E340FFFFFFFFFFFFFFFF",
		x"E35BE35AE359E358E357E356E355E354E353E352E351E350E34FE34EE34DE34C",
		x"E36BE36AE369E368E367E366E365E364E363E362E361E360E35FE35EE35DE35C",
		x"E37BE37AE379E378E377E376E375E374E373E372E371E370E36FE36EE36DE36C",
		x"E387E386E385E384E383E382E381E380FFFFFFFFFFFFFFFFE37FE37EE37DE37C",
		x"E397E396E395E394E393E392E391E390E38FE38EE38DE38CE38BE38AE389E388",
		x"E3A7E3A6E3A5E3A4E3A3E3A2E3A1E3A0E39FE39EE39DE39CE39BE39AE399E398",
		x"E3B7E3B6E3B5E3B4E3B3E3B2E3B1E3B0E3AFE3AEE3ADE3ACE3ABE3AAE3A9E3A8",
		x"E3C3E3C2E3C1E3C0FFFFFFFFFFFFFFFFE3BFE3BEE3BDE3BCE3BBE3BAE3B9E3B8",
		x"E3D3E3D2E3D1E3D0E3CFE3CEE3CDE3CCE3CBE3CAE3C9E3C8E3C7E3C6E3C5E3C4",
		x"E3E3E3E2E3E1E3E0E3DFE3DEE3DDE3DCE3DBE3DAE3D9E3D8E3D7E3D6E3D5E3D4",
		x"E3F3E3F2E3F1E3F0E3EFE3EEE3EDE3ECE3EBE3EAE3E9E3E8E3E7E3E6E3E5E3E4",
		x"FFFFFFFFFFFFFFFFE3FFE3FEE3FDE3FCE3FBE3FAE3F9E3F8E3F7E3F6E3F5E3F4",
		x"E40FE40EE40DE40CE40BE40AE409E408E407E406E405E404E403E402E401E400",
		x"E41FE41EE41DE41CE41BE41AE419E418E417E416E415E414E413E412E411E410",
		x"E42FE42EE42DE42CE42BE42AE429E428E427E426E425E424E423E422E421E420",
		x"E43FE43EE43DE43CE43BE43AE439E438E437E436E435E434E433E432E431E430",
		x"E44BE44AE449E448E447E446E445E444E443E442E441E440FFFFFFFFFFFFFFFF",
		x"E45BE45AE459E458E457E456E455E454E453E452E451E450E44FE44EE44DE44C",
		x"E46BE46AE469E468E467E466E465E464E463E462E461E460E45FE45EE45DE45C",
		x"E47BE47AE479E478E477E476E475E474E473E472E471E470E46FE46EE46DE46C",
		x"E487E486E485E484E483E482E481E480FFFFFFFFFFFFFFFFE47FE47EE47DE47C",
		x"E497E496E495E494E493E492E491E490E48FE48EE48DE48CE48BE48AE489E488",
		x"E4A7E4A6E4A5E4A4E4A3E4A2E4A1E4A0E49FE49EE49DE49CE49BE49AE499E498",
		x"E4B7E4B6E4B5E4B4E4B3E4B2E4B1E4B0E4AFE4AEE4ADE4ACE4ABE4AAE4A9E4A8",
		x"E4C3E4C2E4C1E4C0FFFFFFFFFFFFFFFFE4BFE4BEE4BDE4BCE4BBE4BAE4B9E4B8",
		x"E4D3E4D2E4D1E4D0E4CFE4CEE4CDE4CCE4CBE4CAE4C9E4C8E4C7E4C6E4C5E4C4",
		x"E4E3E4E2E4E1E4E0E4DFE4DEE4DDE4DCE4DBE4DAE4D9E4D8E4D7E4D6E4D5E4D4",
		x"E4F3E4F2E4F1E4F0E4EFE4EEE4EDE4ECE4EBE4EAE4E9E4E8E4E7E4E6E4E5E4E4",
		x"FFFFFFFFFFFFFFFFE4FFE4FEE4FDE4FCE4FBE4FAE4F9E4F8E4F7E4F6E4F5E4F4",
		x"E50FE50EE50DE50CE50BE50AE509E508E507E506E505E504E503E502E501E500",
		x"E51FE51EE51DE51CE51BE51AE519E518E517E516E515E514E513E512E511E510",
		x"E52FE52EE52DE52CE52BE52AE529E528E527E526E525E524E523E522E521E520",
		x"E53FE53EE53DE53CE53BE53AE539E538E537E536E535E534E533E532E531E530",
		x"E54BE54AE549E548E547E546E545E544E543E542E541E540FFFFFFFFFFFFFFFF",
		x"E55BE55AE559E558E557E556E555E554E553E552E551E550E54FE54EE54DE54C",
		x"E56BE56AE569E568E567E566E565E564E563E562E561E560E55FE55EE55DE55C",
		x"E57BE57AE579E578E577E576E575E574E573E572E571E570E56FE56EE56DE56C",
		x"E587E586E585E584E583E582E581E580FFFFFFFFFFFFFFFFE57FE57EE57DE57C",
		x"E597E596E595E594E593E592E591E590E58FE58EE58DE58CE58BE58AE589E588",
		x"E5A7E5A6E5A5E5A4E5A3E5A2E5A1E5A0E59FE59EE59DE59CE59BE59AE599E598",
		x"E5B7E5B6E5B5E5B4E5B3E5B2E5B1E5B0E5AFE5AEE5ADE5ACE5ABE5AAE5A9E5A8",
		x"E5C3E5C2E5C1E5C0FFFFFFFFFFFFFFFFE5BFE5BEE5BDE5BCE5BBE5BAE5B9E5B8",
		x"E5D3E5D2E5D1E5D0E5CFE5CEE5CDE5CCE5CBE5CAE5C9E5C8E5C7E5C6E5C5E5C4",
		x"E5E3E5E2E5E1E5E0E5DFE5DEE5DDE5DCE5DBE5DAE5D9E5D8E5D7E5D6E5D5E5D4",
		x"E5F3E5F2E5F1E5F0E5EFE5EEE5EDE5ECE5EBE5EAE5E9E5E8E5E7E5E6E5E5E5E4",
		x"FFFFFFFFFFFFFFFFE5FFE5FEE5FDE5FCE5FBE5FAE5F9E5F8E5F7E5F6E5F5E5F4",
		x"E60FE60EE60DE60CE60BE60AE609E608E607E606E605E604E603E602E601E600",
		x"E61FE61EE61DE61CE61BE61AE619E618E617E616E615E614E613E612E611E610",
		x"E62FE62EE62DE62CE62BE62AE629E628E627E626E625E624E623E622E621E620",
		x"E63FE63EE63DE63CE63BE63AE639E638E637E636E635E634E633E632E631E630",
		x"E64BE64AE649E648E647E646E645E644E643E642E641E640FFFFFFFFFFFFFFFF",
		x"E65BE65AE659E658E657E656E655E654E653E652E651E650E64FE64EE64DE64C",
		x"E66BE66AE669E668E667E666E665E664E663E662E661E660E65FE65EE65DE65C",
		x"E67BE67AE679E678E677E676E675E674E673E672E671E670E66FE66EE66DE66C",
		x"E687E686E685E684E683E682E681E680FFFFFFFFFFFFFFFFE67FE67EE67DE67C",
		x"E697E696E695E694E693E692E691E690E68FE68EE68DE68CE68BE68AE689E688",
		x"E6A7E6A6E6A5E6A4E6A3E6A2E6A1E6A0E69FE69EE69DE69CE69BE69AE699E698",
		x"E6B7E6B6E6B5E6B4E6B3E6B2E6B1E6B0E6AFE6AEE6ADE6ACE6ABE6AAE6A9E6A8",
		x"E6C3E6C2E6C1E6C0FFFFFFFFFFFFFFFFE6BFE6BEE6BDE6BCE6BBE6BAE6B9E6B8",
		x"E6D3E6D2E6D1E6D0E6CFE6CEE6CDE6CCE6CBE6CAE6C9E6C8E6C7E6C6E6C5E6C4",
		x"E6E3E6E2E6E1E6E0E6DFE6DEE6DDE6DCE6DBE6DAE6D9E6D8E6D7E6D6E6D5E6D4",
		x"E6F3E6F2E6F1E6F0E6EFE6EEE6EDE6ECE6EBE6EAE6E9E6E8E6E7E6E6E6E5E6E4",
		x"FFFFFFFFFFFFFFFFE6FFE6FEE6FDE6FCE6FBE6FAE6F9E6F8E6F7E6F6E6F5E6F4",
		x"E70FE70EE70DE70CE70BE70AE709E708E707E706E705E704E703E702E701E700",
		x"E71FE71EE71DE71CE71BE71AE719E718E717E716E715E714E713E712E711E710",
		x"E72FE72EE72DE72CE72BE72AE729E728E727E726E725E724E723E722E721E720",
		x"E73FE73EE73DE73CE73BE73AE739E738E737E736E735E734E733E732E731E730",
		x"E74BE74AE749E748E747E746E745E744E743E742E741E740FFFFFFFFFFFFFFFF",
		x"E75BE75AE759E758E757E756E755E754E753E752E751E750E74FE74EE74DE74C",
		x"E76BE76AE769E768E767E766E765E764E763E762E761E760E75FE75EE75DE75C",
		x"E77BE77AE779E778E777E776E775E774E773E772E771E770E76FE76EE76DE76C",
		x"E787E786E785E784E783E782E781E780FFFFFFFFFFFFFFFFE77FE77EE77DE77C",
		x"E797E796E795E794E793E792E791E790E78FE78EE78DE78CE78BE78AE789E788",
		x"E7A7E7A6E7A5E7A4E7A3E7A2E7A1E7A0E79FE79EE79DE79CE79BE79AE799E798",
		x"E7B7E7B6E7B5E7B4E7B3E7B2E7B1E7B0E7AFE7AEE7ADE7ACE7ABE7AAE7A9E7A8",
		x"E7C3E7C2E7C1E7C0FFFFFFFFFFFFFFFFE7BFE7BEE7BDE7BCE7BBE7BAE7B9E7B8",
		x"E7D3E7D2E7D1E7D0E7CFE7CEE7CDE7CCE7CBE7CAE7C9E7C8E7C7E7C6E7C5E7C4",
		x"E7E3E7E2E7E1E7E0E7DFE7DEE7DDE7DCE7DBE7DAE7D9E7D8E7D7E7D6E7D5E7D4",
		x"E7F3E7F2E7F1E7F0E7EFE7EEE7EDE7ECE7EBE7EAE7E9E7E8E7E7E7E6E7E5E7E4",
		x"FFFFFFFFFFFFFFFFE7FFE7FEE7FDE7FCE7FBE7FAE7F9E7F8E7F7E7F6E7F5E7F4",
		x"E80FE80EE80DE80CE80BE80AE809E808E807E806E805E804E803E802E801E800",
		x"E81FE81EE81DE81CE81BE81AE819E818E817E816E815E814E813E812E811E810",
		x"E82FE82EE82DE82CE82BE82AE829E828E827E826E825E824E823E822E821E820",
		x"E83FE83EE83DE83CE83BE83AE839E838E837E836E835E834E833E832E831E830",
		x"E84BE84AE849E848E847E846E845E844E843E842E841E840FFFFFFFFFFFFFFFF",
		x"E85BE85AE859E858E857E856E855E854E853E852E851E850E84FE84EE84DE84C",
		x"E86BE86AE869E868E867E866E865E864E863E862E861E860E85FE85EE85DE85C",
		x"E87BE87AE879E878E877E876E875E874E873E872E871E870E86FE86EE86DE86C",
		x"E887E886E885E884E883E882E881E880FFFFFFFFFFFFFFFFE87FE87EE87DE87C",
		x"E897E896E895E894E893E892E891E890E88FE88EE88DE88CE88BE88AE889E888",
		x"E8A7E8A6E8A5E8A4E8A3E8A2E8A1E8A0E89FE89EE89DE89CE89BE89AE899E898",
		x"E8B7E8B6E8B5E8B4E8B3E8B2E8B1E8B0E8AFE8AEE8ADE8ACE8ABE8AAE8A9E8A8",
		x"E8C3E8C2E8C1E8C0FFFFFFFFFFFFFFFFE8BFE8BEE8BDE8BCE8BBE8BAE8B9E8B8",
		x"E8D3E8D2E8D1E8D0E8CFE8CEE8CDE8CCE8CBE8CAE8C9E8C8E8C7E8C6E8C5E8C4",
		x"E8E3E8E2E8E1E8E0E8DFE8DEE8DDE8DCE8DBE8DAE8D9E8D8E8D7E8D6E8D5E8D4",
		x"E8F3E8F2E8F1E8F0E8EFE8EEE8EDE8ECE8EBE8EAE8E9E8E8E8E7E8E6E8E5E8E4",
		x"FFFFFFFFFFFFFFFFE8FFE8FEE8FDE8FCE8FBE8FAE8F9E8F8E8F7E8F6E8F5E8F4",
		x"E90FE90EE90DE90CE90BE90AE909E908E907E906E905E904E903E902E901E900",
		x"E91FE91EE91DE91CE91BE91AE919E918E917E916E915E914E913E912E911E910",
		x"E92FE92EE92DE92CE92BE92AE929E928E927E926E925E924E923E922E921E920",
		x"E93FE93EE93DE93CE93BE93AE939E938E937E936E935E934E933E932E931E930",
		x"E94BE94AE949E948E947E946E945E944E943E942E941E940FFFFFFFFFFFFFFFF",
		x"E95BE95AE959E958E957E956E955E954E953E952E951E950E94FE94EE94DE94C",
		x"E96BE96AE969E968E967E966E965E964E963E962E961E960E95FE95EE95DE95C",
		x"E97BE97AE979E978E977E976E975E974E973E972E971E970E96FE96EE96DE96C",
		x"E987E986E985E984E983E982E981E980FFFFFFFFFFFFFFFFE97FE97EE97DE97C",
		x"E997E996E995E994E993E992E991E990E98FE98EE98DE98CE98BE98AE989E988",
		x"E9A7E9A6E9A5E9A4E9A3E9A2E9A1E9A0E99FE99EE99DE99CE99BE99AE999E998",
		x"E9B7E9B6E9B5E9B4E9B3E9B2E9B1E9B0E9AFE9AEE9ADE9ACE9ABE9AAE9A9E9A8",
		x"E9C3E9C2E9C1E9C0FFFFFFFFFFFFFFFFE9BFE9BEE9BDE9BCE9BBE9BAE9B9E9B8",
		x"E9D3E9D2E9D1E9D0E9CFE9CEE9CDE9CCE9CBE9CAE9C9E9C8E9C7E9C6E9C5E9C4",
		x"E9E3E9E2E9E1E9E0E9DFE9DEE9DDE9DCE9DBE9DAE9D9E9D8E9D7E9D6E9D5E9D4",
		x"E9F3E9F2E9F1E9F0E9EFE9EEE9EDE9ECE9EBE9EAE9E9E9E8E9E7E9E6E9E5E9E4",
		x"FFFFFFFFFFFFFFFFE9FFE9FEE9FDE9FCE9FBE9FAE9F9E9F8E9F7E9F6E9F5E9F4",
		x"EA0FEA0EEA0DEA0CEA0BEA0AEA09EA08EA07EA06EA05EA04EA03EA02EA01EA00",
		x"EA1FEA1EEA1DEA1CEA1BEA1AEA19EA18EA17EA16EA15EA14EA13EA12EA11EA10",
		x"EA2FEA2EEA2DEA2CEA2BEA2AEA29EA28EA27EA26EA25EA24EA23EA22EA21EA20",
		x"EA3FEA3EEA3DEA3CEA3BEA3AEA39EA38EA37EA36EA35EA34EA33EA32EA31EA30",
		x"EA4BEA4AEA49EA48EA47EA46EA45EA44EA43EA42EA41EA40FFFFFFFFFFFFFFFF",
		x"EA5BEA5AEA59EA58EA57EA56EA55EA54EA53EA52EA51EA50EA4FEA4EEA4DEA4C",
		x"EA6BEA6AEA69EA68EA67EA66EA65EA64EA63EA62EA61EA60EA5FEA5EEA5DEA5C",
		x"EA7BEA7AEA79EA78EA77EA76EA75EA74EA73EA72EA71EA70EA6FEA6EEA6DEA6C",
		x"EA87EA86EA85EA84EA83EA82EA81EA80FFFFFFFFFFFFFFFFEA7FEA7EEA7DEA7C",
		x"EA97EA96EA95EA94EA93EA92EA91EA90EA8FEA8EEA8DEA8CEA8BEA8AEA89EA88",
		x"EAA7EAA6EAA5EAA4EAA3EAA2EAA1EAA0EA9FEA9EEA9DEA9CEA9BEA9AEA99EA98",
		x"EAB7EAB6EAB5EAB4EAB3EAB2EAB1EAB0EAAFEAAEEAADEAACEAABEAAAEAA9EAA8",
		x"EAC3EAC2EAC1EAC0FFFFFFFFFFFFFFFFEABFEABEEABDEABCEABBEABAEAB9EAB8",
		x"EAD3EAD2EAD1EAD0EACFEACEEACDEACCEACBEACAEAC9EAC8EAC7EAC6EAC5EAC4",
		x"EAE3EAE2EAE1EAE0EADFEADEEADDEADCEADBEADAEAD9EAD8EAD7EAD6EAD5EAD4",
		x"EAF3EAF2EAF1EAF0EAEFEAEEEAEDEAECEAEBEAEAEAE9EAE8EAE7EAE6EAE5EAE4",
		x"FFFFFFFFFFFFFFFFEAFFEAFEEAFDEAFCEAFBEAFAEAF9EAF8EAF7EAF6EAF5EAF4",
		x"EB0FEB0EEB0DEB0CEB0BEB0AEB09EB08EB07EB06EB05EB04EB03EB02EB01EB00",
		x"EB1FEB1EEB1DEB1CEB1BEB1AEB19EB18EB17EB16EB15EB14EB13EB12EB11EB10",
		x"EB2FEB2EEB2DEB2CEB2BEB2AEB29EB28EB27EB26EB25EB24EB23EB22EB21EB20",
		x"EB3FEB3EEB3DEB3CEB3BEB3AEB39EB38EB37EB36EB35EB34EB33EB32EB31EB30",
		x"EB4BEB4AEB49EB48EB47EB46EB45EB44EB43EB42EB41EB40FFFFFFFFFFFFFFFF",
		x"EB5BEB5AEB59EB58EB57EB56EB55EB54EB53EB52EB51EB50EB4FEB4EEB4DEB4C",
		x"EB6BEB6AEB69EB68EB67EB66EB65EB64EB63EB62EB61EB60EB5FEB5EEB5DEB5C",
		x"EB7BEB7AEB79EB78EB77EB76EB75EB74EB73EB72EB71EB70EB6FEB6EEB6DEB6C",
		x"EB87EB86EB85EB84EB83EB82EB81EB80FFFFFFFFFFFFFFFFEB7FEB7EEB7DEB7C",
		x"EB97EB96EB95EB94EB93EB92EB91EB90EB8FEB8EEB8DEB8CEB8BEB8AEB89EB88",
		x"EBA7EBA6EBA5EBA4EBA3EBA2EBA1EBA0EB9FEB9EEB9DEB9CEB9BEB9AEB99EB98",
		x"EBB7EBB6EBB5EBB4EBB3EBB2EBB1EBB0EBAFEBAEEBADEBACEBABEBAAEBA9EBA8",
		x"EBC3EBC2EBC1EBC0FFFFFFFFFFFFFFFFEBBFEBBEEBBDEBBCEBBBEBBAEBB9EBB8",
		x"EBD3EBD2EBD1EBD0EBCFEBCEEBCDEBCCEBCBEBCAEBC9EBC8EBC7EBC6EBC5EBC4",
		x"EBE3EBE2EBE1EBE0EBDFEBDEEBDDEBDCEBDBEBDAEBD9EBD8EBD7EBD6EBD5EBD4",
		x"EBF3EBF2EBF1EBF0EBEFEBEEEBEDEBECEBEBEBEAEBE9EBE8EBE7EBE6EBE5EBE4",
		x"FFFFFFFFFFFFFFFFEBFFEBFEEBFDEBFCEBFBEBFAEBF9EBF8EBF7EBF6EBF5EBF4",
		x"EC0FEC0EEC0DEC0CEC0BEC0AEC09EC08EC07EC06EC05EC04EC03EC02EC01EC00",
		x"EC1FEC1EEC1DEC1CEC1BEC1AEC19EC18EC17EC16EC15EC14EC13EC12EC11EC10",
		x"EC2FEC2EEC2DEC2CEC2BEC2AEC29EC28EC27EC26EC25EC24EC23EC22EC21EC20",
		x"EC3FEC3EEC3DEC3CEC3BEC3AEC39EC38EC37EC36EC35EC34EC33EC32EC31EC30",
		x"EC4BEC4AEC49EC48EC47EC46EC45EC44EC43EC42EC41EC40FFFFFFFFFFFFFFFF",
		x"EC5BEC5AEC59EC58EC57EC56EC55EC54EC53EC52EC51EC50EC4FEC4EEC4DEC4C",
		x"EC6BEC6AEC69EC68EC67EC66EC65EC64EC63EC62EC61EC60EC5FEC5EEC5DEC5C",
		x"EC7BEC7AEC79EC78EC77EC76EC75EC74EC73EC72EC71EC70EC6FEC6EEC6DEC6C",
		x"EC87EC86EC85EC84EC83EC82EC81EC80FFFFFFFFFFFFFFFFEC7FEC7EEC7DEC7C",
		x"EC97EC96EC95EC94EC93EC92EC91EC90EC8FEC8EEC8DEC8CEC8BEC8AEC89EC88",
		x"ECA7ECA6ECA5ECA4ECA3ECA2ECA1ECA0EC9FEC9EEC9DEC9CEC9BEC9AEC99EC98",
		x"ECB7ECB6ECB5ECB4ECB3ECB2ECB1ECB0ECAFECAEECADECACECABECAAECA9ECA8",
		x"ECC3ECC2ECC1ECC0FFFFFFFFFFFFFFFFECBFECBEECBDECBCECBBECBAECB9ECB8",
		x"ECD3ECD2ECD1ECD0ECCFECCEECCDECCCECCBECCAECC9ECC8ECC7ECC6ECC5ECC4",
		x"ECE3ECE2ECE1ECE0ECDFECDEECDDECDCECDBECDAECD9ECD8ECD7ECD6ECD5ECD4",
		x"ECF3ECF2ECF1ECF0ECEFECEEECEDECECECEBECEAECE9ECE8ECE7ECE6ECE5ECE4",
		x"FFFFFFFFFFFFFFFFECFFECFEECFDECFCECFBECFAECF9ECF8ECF7ECF6ECF5ECF4",
		x"ED0FED0EED0DED0CED0BED0AED09ED08ED07ED06ED05ED04ED03ED02ED01ED00",
		x"ED1FED1EED1DED1CED1BED1AED19ED18ED17ED16ED15ED14ED13ED12ED11ED10",
		x"ED2FED2EED2DED2CED2BED2AED29ED28ED27ED26ED25ED24ED23ED22ED21ED20",
		x"ED3FED3EED3DED3CED3BED3AED39ED38ED37ED36ED35ED34ED33ED32ED31ED30",
		x"ED4BED4AED49ED48ED47ED46ED45ED44ED43ED42ED41ED40FFFFFFFFFFFFFFFF",
		x"ED5BED5AED59ED58ED57ED56ED55ED54ED53ED52ED51ED50ED4FED4EED4DED4C",
		x"ED6BED6AED69ED68ED67ED66ED65ED64ED63ED62ED61ED60ED5FED5EED5DED5C",
		x"ED7BED7AED79ED78ED77ED76ED75ED74ED73ED72ED71ED70ED6FED6EED6DED6C",
		x"ED87ED86ED85ED84ED83ED82ED81ED80FFFFFFFFFFFFFFFFED7FED7EED7DED7C",
		x"ED97ED96ED95ED94ED93ED92ED91ED90ED8FED8EED8DED8CED8BED8AED89ED88",
		x"EDA7EDA6EDA5EDA4EDA3EDA2EDA1EDA0ED9FED9EED9DED9CED9BED9AED99ED98",
		x"EDB7EDB6EDB5EDB4EDB3EDB2EDB1EDB0EDAFEDAEEDADEDACEDABEDAAEDA9EDA8",
		x"EDC3EDC2EDC1EDC0FFFFFFFFFFFFFFFFEDBFEDBEEDBDEDBCEDBBEDBAEDB9EDB8",
		x"EDD3EDD2EDD1EDD0EDCFEDCEEDCDEDCCEDCBEDCAEDC9EDC8EDC7EDC6EDC5EDC4",
		x"EDE3EDE2EDE1EDE0EDDFEDDEEDDDEDDCEDDBEDDAEDD9EDD8EDD7EDD6EDD5EDD4",
		x"EDF3EDF2EDF1EDF0EDEFEDEEEDEDEDECEDEBEDEAEDE9EDE8EDE7EDE6EDE5EDE4",
		x"FFFFFFFFFFFFFFFFEDFFEDFEEDFDEDFCEDFBEDFAEDF9EDF8EDF7EDF6EDF5EDF4",
		x"EE0FEE0EEE0DEE0CEE0BEE0AEE09EE08EE07EE06EE05EE04EE03EE02EE01EE00",
		x"EE1FEE1EEE1DEE1CEE1BEE1AEE19EE18EE17EE16EE15EE14EE13EE12EE11EE10",
		x"EE2FEE2EEE2DEE2CEE2BEE2AEE29EE28EE27EE26EE25EE24EE23EE22EE21EE20",
		x"EE3FEE3EEE3DEE3CEE3BEE3AEE39EE38EE37EE36EE35EE34EE33EE32EE31EE30",
		x"EE4BEE4AEE49EE48EE47EE46EE45EE44EE43EE42EE41EE40FFFFFFFFFFFFFFFF",
		x"EE5BEE5AEE59EE58EE57EE56EE55EE54EE53EE52EE51EE50EE4FEE4EEE4DEE4C",
		x"EE6BEE6AEE69EE68EE67EE66EE65EE64EE63EE62EE61EE60EE5FEE5EEE5DEE5C",
		x"EE7BEE7AEE79EE78EE77EE76EE75EE74EE73EE72EE71EE70EE6FEE6EEE6DEE6C",
		x"EE87EE86EE85EE84EE83EE82EE81EE80FFFFFFFFFFFFFFFFEE7FEE7EEE7DEE7C",
		x"EE97EE96EE95EE94EE93EE92EE91EE90EE8FEE8EEE8DEE8CEE8BEE8AEE89EE88",
		x"EEA7EEA6EEA5EEA4EEA3EEA2EEA1EEA0EE9FEE9EEE9DEE9CEE9BEE9AEE99EE98",
		x"EEB7EEB6EEB5EEB4EEB3EEB2EEB1EEB0EEAFEEAEEEADEEACEEABEEAAEEA9EEA8",
		x"EEC3EEC2EEC1EEC0FFFFFFFFFFFFFFFFEEBFEEBEEEBDEEBCEEBBEEBAEEB9EEB8",
		x"EED3EED2EED1EED0EECFEECEEECDEECCEECBEECAEEC9EEC8EEC7EEC6EEC5EEC4",
		x"EEE3EEE2EEE1EEE0EEDFEEDEEEDDEEDCEEDBEEDAEED9EED8EED7EED6EED5EED4",
		x"EEF3EEF2EEF1EEF0EEEFEEEEEEEDEEECEEEBEEEAEEE9EEE8EEE7EEE6EEE5EEE4",
		x"FFFFFFFFFFFFFFFFEEFFEEFEEEFDEEFCEEFBEEFAEEF9EEF8EEF7EEF6EEF5EEF4",
		x"EF0FEF0EEF0DEF0CEF0BEF0AEF09EF08EF07EF06EF05EF04EF03EF02EF01EF00",
		x"EF1FEF1EEF1DEF1CEF1BEF1AEF19EF18EF17EF16EF15EF14EF13EF12EF11EF10",
		x"EF2FEF2EEF2DEF2CEF2BEF2AEF29EF28EF27EF26EF25EF24EF23EF22EF21EF20",
		x"EF3FEF3EEF3DEF3CEF3BEF3AEF39EF38EF37EF36EF35EF34EF33EF32EF31EF30",
		x"EF4BEF4AEF49EF48EF47EF46EF45EF44EF43EF42EF41EF40FFFFFFFFFFFFFFFF",
		x"EF5BEF5AEF59EF58EF57EF56EF55EF54EF53EF52EF51EF50EF4FEF4EEF4DEF4C",
		x"EF6BEF6AEF69EF68EF67EF66EF65EF64EF63EF62EF61EF60EF5FEF5EEF5DEF5C",
		x"EF7BEF7AEF79EF78EF77EF76EF75EF74EF73EF72EF71EF70EF6FEF6EEF6DEF6C",
		x"EF87EF86EF85EF84EF83EF82EF81EF80FFFFFFFFFFFFFFFFEF7FEF7EEF7DEF7C",
		x"EF97EF96EF95EF94EF93EF92EF91EF90EF8FEF8EEF8DEF8CEF8BEF8AEF89EF88",
		x"EFA7EFA6EFA5EFA4EFA3EFA2EFA1EFA0EF9FEF9EEF9DEF9CEF9BEF9AEF99EF98",
		x"EFB7EFB6EFB5EFB4EFB3EFB2EFB1EFB0EFAFEFAEEFADEFACEFABEFAAEFA9EFA8",
		x"EFC3EFC2EFC1EFC0FFFFFFFFFFFFFFFFEFBFEFBEEFBDEFBCEFBBEFBAEFB9EFB8",
		x"EFD3EFD2EFD1EFD0EFCFEFCEEFCDEFCCEFCBEFCAEFC9EFC8EFC7EFC6EFC5EFC4",
		x"EFE3EFE2EFE1EFE0EFDFEFDEEFDDEFDCEFDBEFDAEFD9EFD8EFD7EFD6EFD5EFD4",
		x"EFF3EFF2EFF1EFF0EFEFEFEEEFEDEFECEFEBEFEAEFE9EFE8EFE7EFE6EFE5EFE4",
		x"FFFFFFFFFFFFFFFFEFFFEFFEEFFDEFFCEFFBEFFAEFF9EFF8EFF7EFF6EFF5EFF4",
		x"F00FF00EF00DF00CF00BF00AF009F008F007F006F005F004F003F002F001F000",
		x"F01FF01EF01DF01CF01BF01AF019F018F017F016F015F014F013F012F011F010",
		x"F02FF02EF02DF02CF02BF02AF029F028F027F026F025F024F023F022F021F020",
		x"F03FF03EF03DF03CF03BF03AF039F038F037F036F035F034F033F032F031F030",
		x"F04BF04AF049F048F047F046F045F044F043F042F041F040FFFFFFFFFFFFFFFF",
		x"F05BF05AF059F058F057F056F055F054F053F052F051F050F04FF04EF04DF04C",
		x"F06BF06AF069F068F067F066F065F064F063F062F061F060F05FF05EF05DF05C",
		x"F07BF07AF079F078F077F076F075F074F073F072F071F070F06FF06EF06DF06C",
		x"F087F086F085F084F083F082F081F080FFFFFFFFFFFFFFFFF07FF07EF07DF07C",
		x"F097F096F095F094F093F092F091F090F08FF08EF08DF08CF08BF08AF089F088",
		x"F0A7F0A6F0A5F0A4F0A3F0A2F0A1F0A0F09FF09EF09DF09CF09BF09AF099F098",
		x"F0B7F0B6F0B5F0B4F0B3F0B2F0B1F0B0F0AFF0AEF0ADF0ACF0ABF0AAF0A9F0A8",
		x"F0C3F0C2F0C1F0C0FFFFFFFFFFFFFFFFF0BFF0BEF0BDF0BCF0BBF0BAF0B9F0B8",
		x"F0D3F0D2F0D1F0D0F0CFF0CEF0CDF0CCF0CBF0CAF0C9F0C8F0C7F0C6F0C5F0C4",
		x"F0E3F0E2F0E1F0E0F0DFF0DEF0DDF0DCF0DBF0DAF0D9F0D8F0D7F0D6F0D5F0D4",
		x"F0F3F0F2F0F1F0F0F0EFF0EEF0EDF0ECF0EBF0EAF0E9F0E8F0E7F0E6F0E5F0E4",
		x"FFFFFFFFFFFFFFFFF0FFF0FEF0FDF0FCF0FBF0FAF0F9F0F8F0F7F0F6F0F5F0F4",
		x"F10FF10EF10DF10CF10BF10AF109F108F107F106F105F104F103F102F101F100",
		x"F11FF11EF11DF11CF11BF11AF119F118F117F116F115F114F113F112F111F110",
		x"F12FF12EF12DF12CF12BF12AF129F128F127F126F125F124F123F122F121F120",
		x"F13FF13EF13DF13CF13BF13AF139F138F137F136F135F134F133F132F131F130",
		x"F14BF14AF149F148F147F146F145F144F143F142F141F140FFFFFFFFFFFFFFFF",
		x"F15BF15AF159F158F157F156F155F154F153F152F151F150F14FF14EF14DF14C",
		x"F16BF16AF169F168F167F166F165F164F163F162F161F160F15FF15EF15DF15C",
		x"F17BF17AF179F178F177F176F175F174F173F172F171F170F16FF16EF16DF16C",
		x"F187F186F185F184F183F182F181F180FFFFFFFFFFFFFFFFF17FF17EF17DF17C",
		x"F197F196F195F194F193F192F191F190F18FF18EF18DF18CF18BF18AF189F188",
		x"F1A7F1A6F1A5F1A4F1A3F1A2F1A1F1A0F19FF19EF19DF19CF19BF19AF199F198",
		x"F1B7F1B6F1B5F1B4F1B3F1B2F1B1F1B0F1AFF1AEF1ADF1ACF1ABF1AAF1A9F1A8",
		x"F1C3F1C2F1C1F1C0FFFFFFFFFFFFFFFFF1BFF1BEF1BDF1BCF1BBF1BAF1B9F1B8",
		x"F1D3F1D2F1D1F1D0F1CFF1CEF1CDF1CCF1CBF1CAF1C9F1C8F1C7F1C6F1C5F1C4",
		x"F1E3F1E2F1E1F1E0F1DFF1DEF1DDF1DCF1DBF1DAF1D9F1D8F1D7F1D6F1D5F1D4",
		x"F1F3F1F2F1F1F1F0F1EFF1EEF1EDF1ECF1EBF1EAF1E9F1E8F1E7F1E6F1E5F1E4",
		x"FFFFFFFFFFFFFFFFF1FFF1FEF1FDF1FCF1FBF1FAF1F9F1F8F1F7F1F6F1F5F1F4",
		x"F20FF20EF20DF20CF20BF20AF209F208F207F206F205F204F203F202F201F200",
		x"F21FF21EF21DF21CF21BF21AF219F218F217F216F215F214F213F212F211F210",
		x"F22FF22EF22DF22CF22BF22AF229F228F227F226F225F224F223F222F221F220",
		x"F23FF23EF23DF23CF23BF23AF239F238F237F236F235F234F233F232F231F230",
		x"F24BF24AF249F248F247F246F245F244F243F242F241F240FFFFFFFFFFFFFFFF",
		x"F25BF25AF259F258F257F256F255F254F253F252F251F250F24FF24EF24DF24C",
		x"F26BF26AF269F268F267F266F265F264F263F262F261F260F25FF25EF25DF25C",
		x"F27BF27AF279F278F277F276F275F274F273F272F271F270F26FF26EF26DF26C",
		x"F287F286F285F284F283F282F281F280FFFFFFFFFFFFFFFFF27FF27EF27DF27C",
		x"F297F296F295F294F293F292F291F290F28FF28EF28DF28CF28BF28AF289F288",
		x"F2A7F2A6F2A5F2A4F2A3F2A2F2A1F2A0F29FF29EF29DF29CF29BF29AF299F298",
		x"F2B7F2B6F2B5F2B4F2B3F2B2F2B1F2B0F2AFF2AEF2ADF2ACF2ABF2AAF2A9F2A8",
		x"F2C3F2C2F2C1F2C0FFFFFFFFFFFFFFFFF2BFF2BEF2BDF2BCF2BBF2BAF2B9F2B8",
		x"F2D3F2D2F2D1F2D0F2CFF2CEF2CDF2CCF2CBF2CAF2C9F2C8F2C7F2C6F2C5F2C4",
		x"F2E3F2E2F2E1F2E0F2DFF2DEF2DDF2DCF2DBF2DAF2D9F2D8F2D7F2D6F2D5F2D4",
		x"F2F3F2F2F2F1F2F0F2EFF2EEF2EDF2ECF2EBF2EAF2E9F2E8F2E7F2E6F2E5F2E4",
		x"FFFFFFFFFFFFFFFFF2FFF2FEF2FDF2FCF2FBF2FAF2F9F2F8F2F7F2F6F2F5F2F4",
		x"F30FF30EF30DF30CF30BF30AF309F308F307F306F305F304F303F302F301F300",
		x"F31FF31EF31DF31CF31BF31AF319F318F317F316F315F314F313F312F311F310",
		x"F32FF32EF32DF32CF32BF32AF329F328F327F326F325F324F323F322F321F320",
		x"F33FF33EF33DF33CF33BF33AF339F338F337F336F335F334F333F332F331F330",
		x"F34BF34AF349F348F347F346F345F344F343F342F341F340FFFFFFFFFFFFFFFF",
		x"F35BF35AF359F358F357F356F355F354F353F352F351F350F34FF34EF34DF34C",
		x"F36BF36AF369F368F367F366F365F364F363F362F361F360F35FF35EF35DF35C",
		x"F37BF37AF379F378F377F376F375F374F373F372F371F370F36FF36EF36DF36C",
		x"F387F386F385F384F383F382F381F380FFFFFFFFFFFFFFFFF37FF37EF37DF37C",
		x"F397F396F395F394F393F392F391F390F38FF38EF38DF38CF38BF38AF389F388",
		x"F3A7F3A6F3A5F3A4F3A3F3A2F3A1F3A0F39FF39EF39DF39CF39BF39AF399F398",
		x"F3B7F3B6F3B5F3B4F3B3F3B2F3B1F3B0F3AFF3AEF3ADF3ACF3ABF3AAF3A9F3A8",
		x"F3C3F3C2F3C1F3C0FFFFFFFFFFFFFFFFF3BFF3BEF3BDF3BCF3BBF3BAF3B9F3B8",
		x"F3D3F3D2F3D1F3D0F3CFF3CEF3CDF3CCF3CBF3CAF3C9F3C8F3C7F3C6F3C5F3C4",
		x"F3E3F3E2F3E1F3E0F3DFF3DEF3DDF3DCF3DBF3DAF3D9F3D8F3D7F3D6F3D5F3D4",
		x"F3F3F3F2F3F1F3F0F3EFF3EEF3EDF3ECF3EBF3EAF3E9F3E8F3E7F3E6F3E5F3E4",
		x"FFFFFFFFFFFFFFFFF3FFF3FEF3FDF3FCF3FBF3FAF3F9F3F8F3F7F3F6F3F5F3F4",
		x"F40FF40EF40DF40CF40BF40AF409F408F407F406F405F404F403F402F401F400",
		x"F41FF41EF41DF41CF41BF41AF419F418F417F416F415F414F413F412F411F410",
		x"F42FF42EF42DF42CF42BF42AF429F428F427F426F425F424F423F422F421F420",
		x"F43FF43EF43DF43CF43BF43AF439F438F437F436F435F434F433F432F431F430",
		x"F44BF44AF449F448F447F446F445F444F443F442F441F440FFFFFFFFFFFFFFFF",
		x"F45BF45AF459F458F457F456F455F454F453F452F451F450F44FF44EF44DF44C",
		x"F46BF46AF469F468F467F466F465F464F463F462F461F460F45FF45EF45DF45C",
		x"F47BF47AF479F478F477F476F475F474F473F472F471F470F46FF46EF46DF46C",
		x"F487F486F485F484F483F482F481F480FFFFFFFFFFFFFFFFF47FF47EF47DF47C",
		x"F497F496F495F494F493F492F491F490F48FF48EF48DF48CF48BF48AF489F488",
		x"F4A7F4A6F4A5F4A4F4A3F4A2F4A1F4A0F49FF49EF49DF49CF49BF49AF499F498",
		x"F4B7F4B6F4B5F4B4F4B3F4B2F4B1F4B0F4AFF4AEF4ADF4ACF4ABF4AAF4A9F4A8",
		x"F4C3F4C2F4C1F4C0FFFFFFFFFFFFFFFFF4BFF4BEF4BDF4BCF4BBF4BAF4B9F4B8",
		x"F4D3F4D2F4D1F4D0F4CFF4CEF4CDF4CCF4CBF4CAF4C9F4C8F4C7F4C6F4C5F4C4",
		x"F4E3F4E2F4E1F4E0F4DFF4DEF4DDF4DCF4DBF4DAF4D9F4D8F4D7F4D6F4D5F4D4",
		x"F4F3F4F2F4F1F4F0F4EFF4EEF4EDF4ECF4EBF4EAF4E9F4E8F4E7F4E6F4E5F4E4",
		x"FFFFFFFFFFFFFFFFF4FFF4FEF4FDF4FCF4FBF4FAF4F9F4F8F4F7F4F6F4F5F4F4",
		x"F50FF50EF50DF50CF50BF50AF509F508F507F506F505F504F503F502F501F500",
		x"F51FF51EF51DF51CF51BF51AF519F518F517F516F515F514F513F512F511F510",
		x"F52FF52EF52DF52CF52BF52AF529F528F527F526F525F524F523F522F521F520",
		x"F53FF53EF53DF53CF53BF53AF539F538F537F536F535F534F533F532F531F530",
		x"F54BF54AF549F548F547F546F545F544F543F542F541F540FFFFFFFFFFFFFFFF",
		x"F55BF55AF559F558F557F556F555F554F553F552F551F550F54FF54EF54DF54C",
		x"F56BF56AF569F568F567F566F565F564F563F562F561F560F55FF55EF55DF55C",
		x"F57BF57AF579F578F577F576F575F574F573F572F571F570F56FF56EF56DF56C",
		x"F587F586F585F584F583F582F581F580FFFFFFFFFFFFFFFFF57FF57EF57DF57C",
		x"F597F596F595F594F593F592F591F590F58FF58EF58DF58CF58BF58AF589F588",
		x"F5A7F5A6F5A5F5A4F5A3F5A2F5A1F5A0F59FF59EF59DF59CF59BF59AF599F598",
		x"F5B7F5B6F5B5F5B4F5B3F5B2F5B1F5B0F5AFF5AEF5ADF5ACF5ABF5AAF5A9F5A8",
		x"F5C3F5C2F5C1F5C0FFFFFFFFFFFFFFFFF5BFF5BEF5BDF5BCF5BBF5BAF5B9F5B8",
		x"F5D3F5D2F5D1F5D0F5CFF5CEF5CDF5CCF5CBF5CAF5C9F5C8F5C7F5C6F5C5F5C4",
		x"F5E3F5E2F5E1F5E0F5DFF5DEF5DDF5DCF5DBF5DAF5D9F5D8F5D7F5D6F5D5F5D4",
		x"F5F3F5F2F5F1F5F0F5EFF5EEF5EDF5ECF5EBF5EAF5E9F5E8F5E7F5E6F5E5F5E4",
		x"FFFFFFFFFFFFFFFFF5FFF5FEF5FDF5FCF5FBF5FAF5F9F5F8F5F7F5F6F5F5F5F4",
		x"F60FF60EF60DF60CF60BF60AF609F608F607F606F605F604F603F602F601F600",
		x"F61FF61EF61DF61CF61BF61AF619F618F617F616F615F614F613F612F611F610",
		x"F62FF62EF62DF62CF62BF62AF629F628F627F626F625F624F623F622F621F620",
		x"F63FF63EF63DF63CF63BF63AF639F638F637F636F635F634F633F632F631F630",
		x"F64BF64AF649F648F647F646F645F644F643F642F641F640FFFFFFFFFFFFFFFF",
		x"F65BF65AF659F658F657F656F655F654F653F652F651F650F64FF64EF64DF64C",
		x"F66BF66AF669F668F667F666F665F664F663F662F661F660F65FF65EF65DF65C",
		x"F67BF67AF679F678F677F676F675F674F673F672F671F670F66FF66EF66DF66C",
		x"F687F686F685F684F683F682F681F680FFFFFFFFFFFFFFFFF67FF67EF67DF67C",
		x"F697F696F695F694F693F692F691F690F68FF68EF68DF68CF68BF68AF689F688",
		x"F6A7F6A6F6A5F6A4F6A3F6A2F6A1F6A0F69FF69EF69DF69CF69BF69AF699F698",
		x"F6B7F6B6F6B5F6B4F6B3F6B2F6B1F6B0F6AFF6AEF6ADF6ACF6ABF6AAF6A9F6A8",
		x"F6C3F6C2F6C1F6C0FFFFFFFFFFFFFFFFF6BFF6BEF6BDF6BCF6BBF6BAF6B9F6B8",
		x"F6D3F6D2F6D1F6D0F6CFF6CEF6CDF6CCF6CBF6CAF6C9F6C8F6C7F6C6F6C5F6C4",
		x"F6E3F6E2F6E1F6E0F6DFF6DEF6DDF6DCF6DBF6DAF6D9F6D8F6D7F6D6F6D5F6D4",
		x"F6F3F6F2F6F1F6F0F6EFF6EEF6EDF6ECF6EBF6EAF6E9F6E8F6E7F6E6F6E5F6E4",
		x"FFFFFFFFFFFFFFFFF6FFF6FEF6FDF6FCF6FBF6FAF6F9F6F8F6F7F6F6F6F5F6F4",
		x"F70FF70EF70DF70CF70BF70AF709F708F707F706F705F704F703F702F701F700",
		x"F71FF71EF71DF71CF71BF71AF719F718F717F716F715F714F713F712F711F710",
		x"F72FF72EF72DF72CF72BF72AF729F728F727F726F725F724F723F722F721F720",
		x"F73FF73EF73DF73CF73BF73AF739F738F737F736F735F734F733F732F731F730",
		x"F74BF74AF749F748F747F746F745F744F743F742F741F740FFFFFFFFFFFFFFFF",
		x"F75BF75AF759F758F757F756F755F754F753F752F751F750F74FF74EF74DF74C",
		x"F76BF76AF769F768F767F766F765F764F763F762F761F760F75FF75EF75DF75C",
		x"F77BF77AF779F778F777F776F775F774F773F772F771F770F76FF76EF76DF76C",
		x"F787F786F785F784F783F782F781F780FFFFFFFFFFFFFFFFF77FF77EF77DF77C",
		x"F797F796F795F794F793F792F791F790F78FF78EF78DF78CF78BF78AF789F788",
		x"F7A7F7A6F7A5F7A4F7A3F7A2F7A1F7A0F79FF79EF79DF79CF79BF79AF799F798",
		x"F7B7F7B6F7B5F7B4F7B3F7B2F7B1F7B0F7AFF7AEF7ADF7ACF7ABF7AAF7A9F7A8",
		x"F7C3F7C2F7C1F7C0FFFFFFFFFFFFFFFFF7BFF7BEF7BDF7BCF7BBF7BAF7B9F7B8",
		x"F7D3F7D2F7D1F7D0F7CFF7CEF7CDF7CCF7CBF7CAF7C9F7C8F7C7F7C6F7C5F7C4",
		x"F7E3F7E2F7E1F7E0F7DFF7DEF7DDF7DCF7DBF7DAF7D9F7D8F7D7F7D6F7D5F7D4",
		x"F7F3F7F2F7F1F7F0F7EFF7EEF7EDF7ECF7EBF7EAF7E9F7E8F7E7F7E6F7E5F7E4",
		x"FFFFFFFFFFFFFFFFF7FFF7FEF7FDF7FCF7FBF7FAF7F9F7F8F7F7F7F6F7F5F7F4",
		x"F80FF80EF80DF80CF80BF80AF809F808F807F806F805F804F803F802F801F800",
		x"F81FF81EF81DF81CF81BF81AF819F818F817F816F815F814F813F812F811F810",
		x"F82FF82EF82DF82CF82BF82AF829F828F827F826F825F824F823F822F821F820",
		x"F83FF83EF83DF83CF83BF83AF839F838F837F836F835F834F833F832F831F830",
		x"F84BF84AF849F848F847F846F845F844F843F842F841F840FFFFFFFFFFFFFFFF",
		x"F85BF85AF859F858F857F856F855F854F853F852F851F850F84FF84EF84DF84C",
		x"F86BF86AF869F868F867F866F865F864F863F862F861F860F85FF85EF85DF85C",
		x"F87BF87AF879F878F877F876F875F874F873F872F871F870F86FF86EF86DF86C",
		x"F887F886F885F884F883F882F881F880FFFFFFFFFFFFFFFFF87FF87EF87DF87C",
		x"F897F896F895F894F893F892F891F890F88FF88EF88DF88CF88BF88AF889F888",
		x"F8A7F8A6F8A5F8A4F8A3F8A2F8A1F8A0F89FF89EF89DF89CF89BF89AF899F898",
		x"F8B7F8B6F8B5F8B4F8B3F8B2F8B1F8B0F8AFF8AEF8ADF8ACF8ABF8AAF8A9F8A8",
		x"F8C3F8C2F8C1F8C0FFFFFFFFFFFFFFFFF8BFF8BEF8BDF8BCF8BBF8BAF8B9F8B8",
		x"F8D3F8D2F8D1F8D0F8CFF8CEF8CDF8CCF8CBF8CAF8C9F8C8F8C7F8C6F8C5F8C4",
		x"F8E3F8E2F8E1F8E0F8DFF8DEF8DDF8DCF8DBF8DAF8D9F8D8F8D7F8D6F8D5F8D4",
		x"F8F3F8F2F8F1F8F0F8EFF8EEF8EDF8ECF8EBF8EAF8E9F8E8F8E7F8E6F8E5F8E4",
		x"FFFFFFFFFFFFFFFFF8FFF8FEF8FDF8FCF8FBF8FAF8F9F8F8F8F7F8F6F8F5F8F4",
		x"F90FF90EF90DF90CF90BF90AF909F908F907F906F905F904F903F902F901F900",
		x"F91FF91EF91DF91CF91BF91AF919F918F917F916F915F914F913F912F911F910",
		x"F92FF92EF92DF92CF92BF92AF929F928F927F926F925F924F923F922F921F920",
		x"F93FF93EF93DF93CF93BF93AF939F938F937F936F935F934F933F932F931F930",
		x"F94BF94AF949F948F947F946F945F944F943F942F941F940FFFFFFFFFFFFFFFF",
		x"F95BF95AF959F958F957F956F955F954F953F952F951F950F94FF94EF94DF94C",
		x"F96BF96AF969F968F967F966F965F964F963F962F961F960F95FF95EF95DF95C",
		x"F97BF97AF979F978F977F976F975F974F973F972F971F970F96FF96EF96DF96C",
		x"F987F986F985F984F983F982F981F980FFFFFFFFFFFFFFFFF97FF97EF97DF97C",
		x"F997F996F995F994F993F992F991F990F98FF98EF98DF98CF98BF98AF989F988",
		x"F9A7F9A6F9A5F9A4F9A3F9A2F9A1F9A0F99FF99EF99DF99CF99BF99AF999F998",
		x"F9B7F9B6F9B5F9B4F9B3F9B2F9B1F9B0F9AFF9AEF9ADF9ACF9ABF9AAF9A9F9A8",
		x"F9C3F9C2F9C1F9C0FFFFFFFFFFFFFFFFF9BFF9BEF9BDF9BCF9BBF9BAF9B9F9B8",
		x"F9D3F9D2F9D1F9D0F9CFF9CEF9CDF9CCF9CBF9CAF9C9F9C8F9C7F9C6F9C5F9C4",
		x"F9E3F9E2F9E1F9E0F9DFF9DEF9DDF9DCF9DBF9DAF9D9F9D8F9D7F9D6F9D5F9D4",
		x"F9F3F9F2F9F1F9F0F9EFF9EEF9EDF9ECF9EBF9EAF9E9F9E8F9E7F9E6F9E5F9E4",
		x"FFFFFFFFFFFFFFFFF9FFF9FEF9FDF9FCF9FBF9FAF9F9F9F8F9F7F9F6F9F5F9F4",
		x"FA0FFA0EFA0DFA0CFA0BFA0AFA09FA08FA07FA06FA05FA04FA03FA02FA01FA00",
		x"FA1FFA1EFA1DFA1CFA1BFA1AFA19FA18FA17FA16FA15FA14FA13FA12FA11FA10",
		x"FA2FFA2EFA2DFA2CFA2BFA2AFA29FA28FA27FA26FA25FA24FA23FA22FA21FA20",
		x"FA3FFA3EFA3DFA3CFA3BFA3AFA39FA38FA37FA36FA35FA34FA33FA32FA31FA30",
		x"FA4BFA4AFA49FA48FA47FA46FA45FA44FA43FA42FA41FA40FFFFFFFFFFFFFFFF",
		x"FA5BFA5AFA59FA58FA57FA56FA55FA54FA53FA52FA51FA50FA4FFA4EFA4DFA4C",
		x"FA6BFA6AFA69FA68FA67FA66FA65FA64FA63FA62FA61FA60FA5FFA5EFA5DFA5C",
		x"FA7BFA7AFA79FA78FA77FA76FA75FA74FA73FA72FA71FA70FA6FFA6EFA6DFA6C",
		x"FA87FA86FA85FA84FA83FA82FA81FA80FFFFFFFFFFFFFFFFFA7FFA7EFA7DFA7C",
		x"FA97FA96FA95FA94FA93FA92FA91FA90FA8FFA8EFA8DFA8CFA8BFA8AFA89FA88",
		x"FAA7FAA6FAA5FAA4FAA3FAA2FAA1FAA0FA9FFA9EFA9DFA9CFA9BFA9AFA99FA98",
		x"FAB7FAB6FAB5FAB4FAB3FAB2FAB1FAB0FAAFFAAEFAADFAACFAABFAAAFAA9FAA8",
		x"FAC3FAC2FAC1FAC0FFFFFFFFFFFFFFFFFABFFABEFABDFABCFABBFABAFAB9FAB8",
		x"FAD3FAD2FAD1FAD0FACFFACEFACDFACCFACBFACAFAC9FAC8FAC7FAC6FAC5FAC4",
		x"FAE3FAE2FAE1FAE0FADFFADEFADDFADCFADBFADAFAD9FAD8FAD7FAD6FAD5FAD4",
		x"FAF3FAF2FAF1FAF0FAEFFAEEFAEDFAECFAEBFAEAFAE9FAE8FAE7FAE6FAE5FAE4",
		x"FFFFFFFFFFFFFFFFFAFFFAFEFAFDFAFCFAFBFAFAFAF9FAF8FAF7FAF6FAF5FAF4",
		x"FB0FFB0EFB0DFB0CFB0BFB0AFB09FB08FB07FB06FB05FB04FB03FB02FB01FB00",
		x"FB1FFB1EFB1DFB1CFB1BFB1AFB19FB18FB17FB16FB15FB14FB13FB12FB11FB10",
		x"FB2FFB2EFB2DFB2CFB2BFB2AFB29FB28FB27FB26FB25FB24FB23FB22FB21FB20",
		x"FB3FFB3EFB3DFB3CFB3BFB3AFB39FB38FB37FB36FB35FB34FB33FB32FB31FB30",
		x"FB4BFB4AFB49FB48FB47FB46FB45FB44FB43FB42FB41FB40FFFFFFFFFFFFFFFF",
		x"FB5BFB5AFB59FB58FB57FB56FB55FB54FB53FB52FB51FB50FB4FFB4EFB4DFB4C",
		x"FB6BFB6AFB69FB68FB67FB66FB65FB64FB63FB62FB61FB60FB5FFB5EFB5DFB5C",
		x"FB7BFB7AFB79FB78FB77FB76FB75FB74FB73FB72FB71FB70FB6FFB6EFB6DFB6C",
		x"FB87FB86FB85FB84FB83FB82FB81FB80FFFFFFFFFFFFFFFFFB7FFB7EFB7DFB7C",
		x"FB97FB96FB95FB94FB93FB92FB91FB90FB8FFB8EFB8DFB8CFB8BFB8AFB89FB88",
		x"FBA7FBA6FBA5FBA4FBA3FBA2FBA1FBA0FB9FFB9EFB9DFB9CFB9BFB9AFB99FB98",
		x"FBB7FBB6FBB5FBB4FBB3FBB2FBB1FBB0FBAFFBAEFBADFBACFBABFBAAFBA9FBA8",
		x"FBC3FBC2FBC1FBC0FFFFFFFFFFFFFFFFFBBFFBBEFBBDFBBCFBBBFBBAFBB9FBB8",
		x"FBD3FBD2FBD1FBD0FBCFFBCEFBCDFBCCFBCBFBCAFBC9FBC8FBC7FBC6FBC5FBC4",
		x"FBE3FBE2FBE1FBE0FBDFFBDEFBDDFBDCFBDBFBDAFBD9FBD8FBD7FBD6FBD5FBD4",
		x"FBF3FBF2FBF1FBF0FBEFFBEEFBEDFBECFBEBFBEAFBE9FBE8FBE7FBE6FBE5FBE4",
		x"FFFFFFFFFFFFFFFFFBFFFBFEFBFDFBFCFBFBFBFAFBF9FBF8FBF7FBF6FBF5FBF4",
		x"FC0FFC0EFC0DFC0CFC0BFC0AFC09FC08FC07FC06FC05FC04FC03FC02FC01FC00",
		x"FC1FFC1EFC1DFC1CFC1BFC1AFC19FC18FC17FC16FC15FC14FC13FC12FC11FC10",
		x"FC2FFC2EFC2DFC2CFC2BFC2AFC29FC28FC27FC26FC25FC24FC23FC22FC21FC20",
		x"FC3FFC3EFC3DFC3CFC3BFC3AFC39FC38FC37FC36FC35FC34FC33FC32FC31FC30",
		x"FC4BFC4AFC49FC48FC47FC46FC45FC44FC43FC42FC41FC40FFFFFFFFFFFFFFFF",
		x"FC5BFC5AFC59FC58FC57FC56FC55FC54FC53FC52FC51FC50FC4FFC4EFC4DFC4C",
		x"FC6BFC6AFC69FC68FC67FC66FC65FC64FC63FC62FC61FC60FC5FFC5EFC5DFC5C",
		x"FC7BFC7AFC79FC78FC77FC76FC75FC74FC73FC72FC71FC70FC6FFC6EFC6DFC6C",
		x"FC87FC86FC85FC84FC83FC82FC81FC80FFFFFFFFFFFFFFFFFC7FFC7EFC7DFC7C",
		x"FC97FC96FC95FC94FC93FC92FC91FC90FC8FFC8EFC8DFC8CFC8BFC8AFC89FC88",
		x"FCA7FCA6FCA5FCA4FCA3FCA2FCA1FCA0FC9FFC9EFC9DFC9CFC9BFC9AFC99FC98",
		x"FCB7FCB6FCB5FCB4FCB3FCB2FCB1FCB0FCAFFCAEFCADFCACFCABFCAAFCA9FCA8",
		x"FCC3FCC2FCC1FCC0FFFFFFFFFFFFFFFFFCBFFCBEFCBDFCBCFCBBFCBAFCB9FCB8",
		x"FCD3FCD2FCD1FCD0FCCFFCCEFCCDFCCCFCCBFCCAFCC9FCC8FCC7FCC6FCC5FCC4",
		x"FCE3FCE2FCE1FCE0FCDFFCDEFCDDFCDCFCDBFCDAFCD9FCD8FCD7FCD6FCD5FCD4",
		x"FCF3FCF2FCF1FCF0FCEFFCEEFCEDFCECFCEBFCEAFCE9FCE8FCE7FCE6FCE5FCE4",
		x"FFFFFFFFFFFFFFFFFCFFFCFEFCFDFCFCFCFBFCFAFCF9FCF8FCF7FCF6FCF5FCF4",
		x"FD0FFD0EFD0DFD0CFD0BFD0AFD09FD08FD07FD06FD05FD04FD03FD02FD01FD00",
		x"FD1FFD1EFD1DFD1CFD1BFD1AFD19FD18FD17FD16FD15FD14FD13FD12FD11FD10",
		x"FD2FFD2EFD2DFD2CFD2BFD2AFD29FD28FD27FD26FD25FD24FD23FD22FD21FD20",
		x"FD3FFD3EFD3DFD3CFD3BFD3AFD39FD38FD37FD36FD35FD34FD33FD32FD31FD30",
		x"FD4BFD4AFD49FD48FD47FD46FD45FD44FD43FD42FD41FD40FFFFFFFFFFFFFFFF",
		x"FD5BFD5AFD59FD58FD57FD56FD55FD54FD53FD52FD51FD50FD4FFD4EFD4DFD4C",
		x"FD6BFD6AFD69FD68FD67FD66FD65FD64FD63FD62FD61FD60FD5FFD5EFD5DFD5C",
		x"FD7BFD7AFD79FD78FD77FD76FD75FD74FD73FD72FD71FD70FD6FFD6EFD6DFD6C",
		x"FD87FD86FD85FD84FD83FD82FD81FD80FFFFFFFFFFFFFFFFFD7FFD7EFD7DFD7C",
		x"FD97FD96FD95FD94FD93FD92FD91FD90FD8FFD8EFD8DFD8CFD8BFD8AFD89FD88",
		x"FDA7FDA6FDA5FDA4FDA3FDA2FDA1FDA0FD9FFD9EFD9DFD9CFD9BFD9AFD99FD98",
		x"FDB7FDB6FDB5FDB4FDB3FDB2FDB1FDB0FDAFFDAEFDADFDACFDABFDAAFDA9FDA8",
		x"FDC3FDC2FDC1FDC0FFFFFFFFFFFFFFFFFDBFFDBEFDBDFDBCFDBBFDBAFDB9FDB8",
		x"FDD3FDD2FDD1FDD0FDCFFDCEFDCDFDCCFDCBFDCAFDC9FDC8FDC7FDC6FDC5FDC4",
		x"FDE3FDE2FDE1FDE0FDDFFDDEFDDDFDDCFDDBFDDAFDD9FDD8FDD7FDD6FDD5FDD4",
		x"FDF3FDF2FDF1FDF0FDEFFDEEFDEDFDECFDEBFDEAFDE9FDE8FDE7FDE6FDE5FDE4",
		x"FFFFFFFFFFFFFFFFFDFFFDFEFDFDFDFCFDFBFDFAFDF9FDF8FDF7FDF6FDF5FDF4",
		x"FE0FFE0EFE0DFE0CFE0BFE0AFE09FE08FE07FE06FE05FE04FE03FE02FE01FE00",
		x"FE1FFE1EFE1DFE1CFE1BFE1AFE19FE18FE17FE16FE15FE14FE13FE12FE11FE10",
		x"FE2FFE2EFE2DFE2CFE2BFE2AFE29FE28FE27FE26FE25FE24FE23FE22FE21FE20",
		x"FE3FFE3EFE3DFE3CFE3BFE3AFE39FE38FE37FE36FE35FE34FE33FE32FE31FE30",
		x"FE4BFE4AFE49FE48FE47FE46FE45FE44FE43FE42FE41FE40FFFFFFFFFFFFFFFF",
		x"FE5BFE5AFE59FE58FE57FE56FE55FE54FE53FE52FE51FE50FE4FFE4EFE4DFE4C",
		x"FE6BFE6AFE69FE68FE67FE66FE65FE64FE63FE62FE61FE60FE5FFE5EFE5DFE5C",
		x"FE7BFE7AFE79FE78FE77FE76FE75FE74FE73FE72FE71FE70FE6FFE6EFE6DFE6C",
		x"FE87FE86FE85FE84FE83FE82FE81FE80FFFFFFFFFFFFFFFFFE7FFE7EFE7DFE7C",
		x"FE97FE96FE95FE94FE93FE92FE91FE90FE8FFE8EFE8DFE8CFE8BFE8AFE89FE88",
		x"FEA7FEA6FEA5FEA4FEA3FEA2FEA1FEA0FE9FFE9EFE9DFE9CFE9BFE9AFE99FE98",
		x"FEB7FEB6FEB5FEB4FEB3FEB2FEB1FEB0FEAFFEAEFEADFEACFEABFEAAFEA9FEA8",
		x"FEC3FEC2FEC1FEC0FFFFFFFFFFFFFFFFFEBFFEBEFEBDFEBCFEBBFEBAFEB9FEB8",
		x"FED3FED2FED1FED0FECFFECEFECDFECCFECBFECAFEC9FEC8FEC7FEC6FEC5FEC4",
		x"FEE3FEE2FEE1FEE0FEDFFEDEFEDDFEDCFEDBFEDAFED9FED8FED7FED6FED5FED4",
		x"FEF3FEF2FEF1FEF0FEEFFEEEFEEDFEECFEEBFEEAFEE9FEE8FEE7FEE6FEE5FEE4",
		x"FFFFFFFFFFFFFFFFFEFFFEFEFEFDFEFCFEFBFEFAFEF9FEF8FEF7FEF6FEF5FEF4",
		x"FF0FFF0EFF0DFF0CFF0BFF0AFF09FF08FF07FF06FF05FF04FF03FF02FF01FF00",
		x"FF1FFF1EFF1DFF1CFF1BFF1AFF19FF18FF17FF16FF15FF14FF13FF12FF11FF10",
		x"FF2FFF2EFF2DFF2CFF2BFF2AFF29FF28FF27FF26FF25FF24FF23FF22FF21FF20",
		x"FF3FFF3EFF3DFF3CFF3BFF3AFF39FF38FF37FF36FF35FF34FF33FF32FF31FF30",
		x"FF4BFF4AFF49FF48FF47FF46FF45FF44FF43FF42FF41FF40FFFFFFFFFFFFFFFF",
		x"FF5BFF5AFF59FF58FF57FF56FF55FF54FF53FF52FF51FF50FF4FFF4EFF4DFF4C",
		x"FF6BFF6AFF69FF68FF67FF66FF65FF64FF63FF62FF61FF60FF5FFF5EFF5DFF5C",
		x"FF7BFF7AFF79FF78FF77FF76FF75FF74FF73FF72FF71FF70FF6FFF6EFF6DFF6C",
		x"FF87FF86FF85FF84FF83FF82FF81FF80FFFFFFFFFFFFFFFFFF7FFF7EFF7DFF7C",
		x"FF97FF96FF95FF94FF93FF92FF91FF90FF8FFF8EFF8DFF8CFF8BFF8AFF89FF88",
		x"FFA7FFA6FFA5FFA4FFA3FFA2FFA1FFA0FF9FFF9EFF9DFF9CFF9BFF9AFF99FF98",
		x"FFB7FFB6FFB5FFB4FFB3FFB2FFB1FFB0FFAFFFAEFFADFFACFFABFFAAFFA9FFA8",
		x"FFC3FFC2FFC1FFC0FFFFFFFFFFFFFFFFFFBFFFBEFFBDFFBCFFBBFFBAFFB9FFB8",
		x"FFD3FFD2FFD1FFD0FFCFFFCEFFCDFFCCFFCBFFCAFFC9FFC8FFC7FFC6FFC5FFC4",
		x"FFE3FFE2FFE1FFE0FFDFFFDEFFDDFFDCFFDBFFDAFFD9FFD8FFD7FFD6FFD5FFD4",
		x"FFF3FFF2FFF1FFF0FFEFFFEEFFEDFFECFFEBFFEAFFE9FFE8FFE7FFE6FFE5FFE4",
		x"FFFFFFFFFFFFFFFFFFFFFFFEFFFDFFFCFFFBFFFAFFF9FFF8FFF7FFF6FFF5FFF4"
	);

	signal s_counter     : natural                                     := 0;
	signal s_address_cnt : natural range 0 to (2**g_ADDRESS_WIDTH - 1) := 0;
	signal s_times_cnt   : natural                                     := 0;

begin

	p_avalon_buffer_R_stimuli : process(clk_i, rst_i) is
	begin
		if (rst_i = '1') then

			avalon_mm_address_o   <= (others => '0');
			avalon_mm_write_o     <= '0';
			avalon_mm_writedata_o <= (others => '0');
			s_ccd_imgdata_cnt     <= 0;
			s_counter             <= 0;
			--						s_counter              <= 5000;
			s_address_cnt         <= 0;
			--			s_mask_cnt             <= 0;
			s_times_cnt           <= 0;

		elsif rising_edge(clk_i) then

			avalon_mm_address_o   <= (others => '0');
			avalon_mm_write_o     <= '0';
			avalon_mm_writedata_o <= (others => '0');
			s_counter             <= s_counter + 1;

			case (s_counter) is

				when 1500 =>
					-- register write
					avalon_mm_address_o   <= std_logic_vector(to_unsigned(s_address_cnt, g_ADDRESS_WIDTH));
					avalon_mm_write_o     <= '1';
					avalon_mm_writedata_o <= c_CCD_IMGDATA(s_ccd_imgdata_cnt);

				when 1501 =>
					if (avalon_mm_waitrequest_i = '1') then
						s_counter <= 1501;
					end if;
					-- register write
					avalon_mm_address_o   <= std_logic_vector(to_unsigned(s_address_cnt, g_ADDRESS_WIDTH));
					avalon_mm_write_o     <= '1';
					avalon_mm_writedata_o <= c_CCD_IMGDATA(s_ccd_imgdata_cnt);

				when 1502 =>
					s_counter     <= 1500;
					if (s_ccd_imgdata_cnt = (c_CCD_IMGDATA_LENGTH - 1)) then
						s_ccd_imgdata_cnt <= 0;
					else
						s_ccd_imgdata_cnt <= s_ccd_imgdata_cnt + 1;
					end if;
					s_address_cnt <= s_address_cnt + 1;
					--if (s_address_cnt = (2**g_ADDRESS_WIDTH - 2)) then
					--					if (s_address_cnt = (1020 - 1)) then
					--					if (s_address_cnt = (272 - 1)) then
					if (s_address_cnt = ((2 ** g_ADDRESS_WIDTH) - 1)) then
						if (s_times_cnt < 1000) then
							s_counter     <= 1500;
							--							s_counter     <= 1000;
							--							s_counter     <= 1500;
							s_address_cnt <= 0;
							s_times_cnt   <= s_times_cnt + 1;
						else
							s_counter     <= 5000;
							s_address_cnt <= 0;
							s_times_cnt   <= 0;
						end if;
					end if;
				--					
				--					if (s_address_cnt = 50) then
				--						s_counter     <= 5000;
				--					end if;

				--				when 1500 =>
				--					-- register write
				--					avalon_mm_address_o   <= std_logic_vector(to_unsigned(s_address_cnt, g_ADDRESS_WIDTH));
				--					avalon_mm_write_o     <= '1';
				--					for cnt in 0 to 3 loop
				--						v_registered_data                                           := (others => '0');
				--						--						if (s_mask_cnt < 16) then
				--						--							s_mask_cnt                      <= s_mask_cnt + 1;
				--						if (v_mask_cnt < 16) then
				--							v_mask_cnt                      := v_mask_cnt + 1;
				--							--						v_registered_data(7 downto 0)   := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							--						v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 2, '1');
				--							--						v_registered_data(15 downto 8)  := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							--						v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 2, '1');
				--							--						v_registered_data(23 downto 16) := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							--						v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 2, '1');
				--							--						v_registered_data(31 downto 24) := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							--						v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 2, '1');
				--							--						v_registered_data(39 downto 32) := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							--						v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 2, '1');
				--							--						v_registered_data(47 downto 40) := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							--						v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 2, '1');
				--							--						v_registered_data(55 downto 48) := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							--						v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 2, '1');
				--							--						v_registered_data(63 downto 56) := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							--						v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 2, '1');
				--							v_registered_data(7 downto 0)   := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 1, '1');
				--							v_registered_data(15 downto 8)  := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 1, '1');
				--							v_registered_data(23 downto 16) := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 1, '1');
				--							v_registered_data(31 downto 24) := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 1, '1');
				--							v_registered_data(39 downto 32) := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 1, '1');
				--							v_registered_data(47 downto 40) := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 1, '1');
				--							v_registered_data(55 downto 48) := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 1, '1');
				--							v_registered_data(63 downto 56) := std_logic_vector(to_unsigned(v_data_cnt, 8));
				--							v_data_cnt                      := f_next_data(v_data_cnt, c_RESET_DATA, c_FINAL_DATA, 1, '1');
				--						else
				--							--							s_mask_cnt        <= 0;
				--							v_mask_cnt        := 0;
				--							--v_registered_data := (others => '1');
				--							--						v_registered_data := x"5555555555555555";
				--							v_registered_data := x"FFFFFFFFFFFFFFFF";
				--						end if;
				--						v_registered_writedata(((64 * cnt) + 63) downto (64 * cnt)) := v_registered_data;
				--					end loop;
				--					avalon_mm_writedata_o <= v_registered_writedata;
				--
				--				when 1501 =>
				--					avalon_mm_address_o   <= std_logic_vector(to_unsigned(s_address_cnt, g_ADDRESS_WIDTH));
				--					avalon_mm_write_o     <= '1';
				--					avalon_mm_writedata_o <= v_registered_writedata;
				--
				--				when 1502 =>
				--					s_counter     <= 1500;
				--					s_address_cnt <= s_address_cnt + 1;
				--					--if (s_address_cnt = (2**g_ADDRESS_WIDTH - 2)) then
				--					--					if (s_address_cnt = (1020 - 1)) then
				--					--					if (s_address_cnt = (272 - 1)) then
				--					if (s_address_cnt = (68 - 1)) then
				----					if (s_address_cnt = (68 - 1)) then
				--						if (s_times_cnt < 1000) then
				--							s_counter     <= 500;
				----							s_counter     <= 1000;
				----							s_counter     <= 1500;
				--							s_address_cnt <= 0;
				--							s_times_cnt   <= s_times_cnt + 1;
				--						else
				--							s_counter     <= 5000;
				--							s_address_cnt <= 0;
				--							s_times_cnt   <= 0;
				--						end if;
				--					end if;

				when others =>
					null;

			end case;

		end if;
	end process p_avalon_buffer_R_stimuli;

end architecture RTL;
