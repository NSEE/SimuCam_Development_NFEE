package rmap_target_write_command_data_eop is
	
end package rmap_target_write_command_data_eop;

package body rmap_target_write_command_data_eop is
	
end package body rmap_target_write_command_data_eop;
