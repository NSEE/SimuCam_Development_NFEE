package rmap_target_write_reply_header_reply_spw_address_pkg is
	
end package rmap_target_write_reply_header_reply_spw_address_pkg;

package body rmap_target_write_reply_header_reply_spw_address_pkg is
	
end package body rmap_target_write_reply_header_reply_spw_address_pkg;
