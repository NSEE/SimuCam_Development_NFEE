// DE4_SOPC.v

// Generated using ACDS version 11.1sp1 216 at 2012.02.03.13:45:47

`timescale 1 ps / 1 ps
module DE4_SOPC (
		output wire        pll_peripheral_clk,                //                         c1_out_clk.clk
		input  wire        reset_n,                           //               ext_clk_clk_in_reset.reset_n
		input  wire [7:0]  in_port_to_the_sw_pio,             //         sw_pio_external_connection.export
		output wire [15:0] out_port_from_the_seven_seg_pio,   //  seven_seg_pio_external_connection.export
		output wire        altpll_0_phasedone_conduit_export, //         altpll_0_phasedone_conduit.export
		output wire [24:0] flash_tristate_bridge_address,     // flash_tristate_bridge_bridge_0_out.flash_tristate_bridge_address
		output wire        flash_tristate_bridge_writen,      //                                   .flash_tristate_bridge_writen
		inout  wire [15:0] flash_tristate_bridge_data,        //                                   .flash_tristate_bridge_data
		output wire        select_n_to_the_ext_flash,         //                                   .select_n_to_the_ext_flash
		output wire        flash_tristate_bridge_readn,       //                                   .flash_tristate_bridge_readn
		output wire        pll_sys_clk,                       //                         c0_out_clk.clk
		input  wire        altpll_0_areset_conduit_export,    //            altpll_0_areset_conduit.export
		output wire        altpll_0_locked_conduit_export,    //            altpll_0_locked_conduit.export
		output wire [7:0]  out_port_from_the_led_pio,         //        led_pio_external_connection.export
		input  wire        ext_clk,                           //                     ext_clk_clk_in.clk
		output wire        mdio_out_from_the_tse_mac,         //         tse_mac_conduit_connection.mdio_out
		output wire        mdio_oen_from_the_tse_mac,         //                                   .mdio_oen
		input  wire        mdio_in_to_the_tse_mac,            //                                   .mdio_in
		output wire        mdc_from_the_tse_mac,              //                                   .mdc
		output wire        led_an_from_the_tse_mac,           //                                   .led_an
		output wire        led_char_err_from_the_tse_mac,     //                                   .led_char_err
		output wire        led_link_from_the_tse_mac,         //                                   .led_link
		output wire        led_disp_err_from_the_tse_mac,     //                                   .led_disp_err
		output wire        led_crs_from_the_tse_mac,          //                                   .led_crs
		output wire        led_col_from_the_tse_mac,          //                                   .led_col
		output wire        txp_from_the_tse_mac,              //                                   .txp
		input  wire        rxp_to_the_tse_mac,                //                                   .rxp
		input  wire        ref_clk_to_the_tse_mac,            //                                   .ref_clk
		output wire        rx_recovclkout_from_the_tse_mac,   //                                   .rx_recovclkout
		input  wire [3:0]  in_port_to_the_pb_pio              //         pb_pio_external_connection.export
	);

	wire         sgdma_tx_out_endofpacket;                                                                          // sgdma_tx:out_endofpacket -> tse_mac:ff_tx_eop
	wire         sgdma_tx_out_valid;                                                                                // sgdma_tx:out_valid -> tse_mac:ff_tx_wren
	wire         sgdma_tx_out_startofpacket;                                                                        // sgdma_tx:out_startofpacket -> tse_mac:ff_tx_sop
	wire         sgdma_tx_out_error;                                                                                // sgdma_tx:out_error -> tse_mac:ff_tx_err
	wire   [1:0] sgdma_tx_out_empty;                                                                                // sgdma_tx:out_empty -> tse_mac:ff_tx_mod
	wire  [31:0] sgdma_tx_out_data;                                                                                 // sgdma_tx:out_data -> tse_mac:ff_tx_data
	wire         sgdma_tx_out_ready;                                                                                // tse_mac:ff_tx_rdy -> sgdma_tx:out_ready
	wire         tse_mac_receive_endofpacket;                                                                       // tse_mac:ff_rx_eop -> sgdma_rx:in_endofpacket
	wire         tse_mac_receive_valid;                                                                             // tse_mac:ff_rx_dval -> sgdma_rx:in_valid
	wire         tse_mac_receive_startofpacket;                                                                     // tse_mac:ff_rx_sop -> sgdma_rx:in_startofpacket
	wire   [5:0] tse_mac_receive_error;                                                                             // tse_mac:rx_err -> sgdma_rx:in_error
	wire   [1:0] tse_mac_receive_empty;                                                                             // tse_mac:ff_rx_mod -> sgdma_rx:in_empty
	wire  [31:0] tse_mac_receive_data;                                                                              // tse_mac:ff_rx_data -> sgdma_rx:in_data
	wire         tse_mac_receive_ready;                                                                             // sgdma_rx:in_ready -> tse_mac:ff_rx_rdy
	wire   [0:0] flash_tristate_bridge_pinsharer_0_tcm_select_n_to_the_ext_flash_out;                               // flash_tristate_bridge_pinSharer_0:select_n_to_the_ext_flash -> flash_tristate_bridge_bridge_0:tcs_select_n_to_the_ext_flash
	wire   [0:0] flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_writen_out;                            // flash_tristate_bridge_pinSharer_0:flash_tristate_bridge_writen -> flash_tristate_bridge_bridge_0:tcs_flash_tristate_bridge_writen
	wire         flash_tristate_bridge_pinsharer_0_tcm_grant;                                                       // flash_tristate_bridge_bridge_0:grant -> flash_tristate_bridge_pinSharer_0:grant
	wire   [0:0] flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_readn_out;                             // flash_tristate_bridge_pinSharer_0:flash_tristate_bridge_readn -> flash_tristate_bridge_bridge_0:tcs_flash_tristate_bridge_readn
	wire  [15:0] flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_out;                              // flash_tristate_bridge_pinSharer_0:flash_tristate_bridge_data -> flash_tristate_bridge_bridge_0:tcs_flash_tristate_bridge_data
	wire         flash_tristate_bridge_pinsharer_0_tcm_request;                                                     // flash_tristate_bridge_pinSharer_0:request -> flash_tristate_bridge_bridge_0:request
	wire         flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_outen;                            // flash_tristate_bridge_pinSharer_0:flash_tristate_bridge_data_outen -> flash_tristate_bridge_bridge_0:tcs_flash_tristate_bridge_data_outen
	wire  [15:0] flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_in;                               // flash_tristate_bridge_bridge_0:tcs_flash_tristate_bridge_data_in -> flash_tristate_bridge_pinSharer_0:flash_tristate_bridge_data_in
	wire  [24:0] flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_address_out;                           // flash_tristate_bridge_pinSharer_0:flash_tristate_bridge_address -> flash_tristate_bridge_bridge_0:tcs_flash_tristate_bridge_address
	wire         ext_flash_tcm_chipselect_n_out;                                                                    // ext_flash:tcm_chipselect_n_out -> flash_tristate_bridge_pinSharer_0:tcs0_chipselect_n_out
	wire         ext_flash_tcm_grant;                                                                               // flash_tristate_bridge_pinSharer_0:tcs0_grant -> ext_flash:tcm_grant
	wire         ext_flash_tcm_data_outen;                                                                          // ext_flash:tcm_data_outen -> flash_tristate_bridge_pinSharer_0:tcs0_data_outen
	wire         ext_flash_tcm_request;                                                                             // ext_flash:tcm_request -> flash_tristate_bridge_pinSharer_0:tcs0_request
	wire  [15:0] ext_flash_tcm_data_out;                                                                            // ext_flash:tcm_data_out -> flash_tristate_bridge_pinSharer_0:tcs0_data_out
	wire         ext_flash_tcm_write_n_out;                                                                         // ext_flash:tcm_write_n_out -> flash_tristate_bridge_pinSharer_0:tcs0_write_n_out
	wire  [24:0] ext_flash_tcm_address_out;                                                                         // ext_flash:tcm_address_out -> flash_tristate_bridge_pinSharer_0:tcs0_address_out
	wire  [15:0] ext_flash_tcm_data_in;                                                                             // flash_tristate_bridge_pinSharer_0:tcs0_data_in -> ext_flash:tcm_data_in
	wire         ext_flash_tcm_read_n_out;                                                                          // ext_flash:tcm_read_n_out -> flash_tristate_bridge_pinSharer_0:tcs0_read_n_out
	wire         cpu_instruction_master_waitrequest;                                                                // cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                                                                    // cpu:i_address -> cpu_instruction_master_translator:av_address
	wire         cpu_instruction_master_read;                                                                       // cpu:i_read -> cpu_instruction_master_translator:av_read
	wire  [31:0] cpu_instruction_master_readdata;                                                                   // cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_readdatavalid;                                                              // cpu_instruction_master_translator:av_readdatavalid -> cpu:i_readdatavalid
	wire         cpu_data_master_waitrequest;                                                                       // cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                                                         // cpu:d_writedata -> cpu_data_master_translator:av_writedata
	wire  [26:0] cpu_data_master_address;                                                                           // cpu:d_address -> cpu_data_master_translator:av_address
	wire         cpu_data_master_write;                                                                             // cpu:d_write -> cpu_data_master_translator:av_write
	wire         cpu_data_master_read;                                                                              // cpu:d_read -> cpu_data_master_translator:av_read
	wire  [31:0] cpu_data_master_readdata;                                                                          // cpu_data_master_translator:av_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                                                                       // cpu:jtag_debug_module_debugaccess_to_roms -> cpu_data_master_translator:av_debugaccess
	wire         cpu_data_master_readdatavalid;                                                                     // cpu_data_master_translator:av_readdatavalid -> cpu:d_readdatavalid
	wire   [3:0] cpu_data_master_byteenable;                                                                        // cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	wire         sgdma_rx_descriptor_read_waitrequest;                                                              // sgdma_rx_descriptor_read_translator:av_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	wire  [31:0] sgdma_rx_descriptor_read_address;                                                                  // sgdma_rx:descriptor_read_address -> sgdma_rx_descriptor_read_translator:av_address
	wire         sgdma_rx_descriptor_read_read;                                                                     // sgdma_rx:descriptor_read_read -> sgdma_rx_descriptor_read_translator:av_read
	wire  [31:0] sgdma_rx_descriptor_read_readdata;                                                                 // sgdma_rx_descriptor_read_translator:av_readdata -> sgdma_rx:descriptor_read_readdata
	wire         sgdma_rx_descriptor_read_readdatavalid;                                                            // sgdma_rx_descriptor_read_translator:av_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	wire         sgdma_rx_descriptor_write_waitrequest;                                                             // sgdma_rx_descriptor_write_translator:av_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	wire  [31:0] sgdma_rx_descriptor_write_writedata;                                                               // sgdma_rx:descriptor_write_writedata -> sgdma_rx_descriptor_write_translator:av_writedata
	wire  [31:0] sgdma_rx_descriptor_write_address;                                                                 // sgdma_rx:descriptor_write_address -> sgdma_rx_descriptor_write_translator:av_address
	wire         sgdma_rx_descriptor_write_write;                                                                   // sgdma_rx:descriptor_write_write -> sgdma_rx_descriptor_write_translator:av_write
	wire         sgdma_tx_descriptor_read_waitrequest;                                                              // sgdma_tx_descriptor_read_translator:av_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	wire  [31:0] sgdma_tx_descriptor_read_address;                                                                  // sgdma_tx:descriptor_read_address -> sgdma_tx_descriptor_read_translator:av_address
	wire         sgdma_tx_descriptor_read_read;                                                                     // sgdma_tx:descriptor_read_read -> sgdma_tx_descriptor_read_translator:av_read
	wire  [31:0] sgdma_tx_descriptor_read_readdata;                                                                 // sgdma_tx_descriptor_read_translator:av_readdata -> sgdma_tx:descriptor_read_readdata
	wire         sgdma_tx_descriptor_read_readdatavalid;                                                            // sgdma_tx_descriptor_read_translator:av_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	wire         sgdma_tx_descriptor_write_waitrequest;                                                             // sgdma_tx_descriptor_write_translator:av_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	wire  [31:0] sgdma_tx_descriptor_write_writedata;                                                               // sgdma_tx:descriptor_write_writedata -> sgdma_tx_descriptor_write_translator:av_writedata
	wire  [31:0] sgdma_tx_descriptor_write_address;                                                                 // sgdma_tx:descriptor_write_address -> sgdma_tx_descriptor_write_translator:av_address
	wire         sgdma_tx_descriptor_write_write;                                                                   // sgdma_tx:descriptor_write_write -> sgdma_tx_descriptor_write_translator:av_write
	wire         sgdma_rx_m_write_waitrequest;                                                                      // sgdma_rx_m_write_translator:av_waitrequest -> sgdma_rx:m_write_waitrequest
	wire  [31:0] sgdma_rx_m_write_writedata;                                                                        // sgdma_rx:m_write_writedata -> sgdma_rx_m_write_translator:av_writedata
	wire  [31:0] sgdma_rx_m_write_address;                                                                          // sgdma_rx:m_write_address -> sgdma_rx_m_write_translator:av_address
	wire         sgdma_rx_m_write_write;                                                                            // sgdma_rx:m_write_write -> sgdma_rx_m_write_translator:av_write
	wire   [3:0] sgdma_rx_m_write_byteenable;                                                                       // sgdma_rx:m_write_byteenable -> sgdma_rx_m_write_translator:av_byteenable
	wire         sgdma_tx_m_read_waitrequest;                                                                       // sgdma_tx_m_read_translator:av_waitrequest -> sgdma_tx:m_read_waitrequest
	wire  [31:0] sgdma_tx_m_read_address;                                                                           // sgdma_tx:m_read_address -> sgdma_tx_m_read_translator:av_address
	wire         sgdma_tx_m_read_read;                                                                              // sgdma_tx:m_read_read -> sgdma_tx_m_read_translator:av_read
	wire  [31:0] sgdma_tx_m_read_readdata;                                                                          // sgdma_tx_m_read_translator:av_readdata -> sgdma_tx:m_read_readdata
	wire         sgdma_tx_m_read_readdatavalid;                                                                     // sgdma_tx_m_read_translator:av_readdatavalid -> sgdma_tx:m_read_readdatavalid
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                    // cpu_jtag_debug_module_translator:av_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                      // cpu_jtag_debug_module_translator:av_address -> cpu:jtag_debug_module_address
	wire         cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                   // cpu_jtag_debug_module_translator:av_chipselect -> cpu:jtag_debug_module_select
	wire         cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                        // cpu_jtag_debug_module_translator:av_write -> cpu:jtag_debug_module_write
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                     // cpu:jtag_debug_module_readdata -> cpu_jtag_debug_module_translator:av_readdata
	wire         cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                // cpu_jtag_debug_module_translator:av_begintransfer -> cpu:jtag_debug_module_begintransfer
	wire         cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                  // cpu_jtag_debug_module_translator:av_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                   // cpu_jtag_debug_module_translator:av_byteenable -> cpu:jtag_debug_module_byteenable
	wire  [31:0] onchip_memory_s1_translator_avalon_anti_slave_0_writedata;                                         // onchip_memory_s1_translator:av_writedata -> onchip_memory:writedata
	wire  [16:0] onchip_memory_s1_translator_avalon_anti_slave_0_address;                                           // onchip_memory_s1_translator:av_address -> onchip_memory:address
	wire         onchip_memory_s1_translator_avalon_anti_slave_0_chipselect;                                        // onchip_memory_s1_translator:av_chipselect -> onchip_memory:chipselect
	wire         onchip_memory_s1_translator_avalon_anti_slave_0_clken;                                             // onchip_memory_s1_translator:av_clken -> onchip_memory:clken
	wire         onchip_memory_s1_translator_avalon_anti_slave_0_write;                                             // onchip_memory_s1_translator:av_write -> onchip_memory:write
	wire  [31:0] onchip_memory_s1_translator_avalon_anti_slave_0_readdata;                                          // onchip_memory:readdata -> onchip_memory_s1_translator:av_readdata
	wire   [3:0] onchip_memory_s1_translator_avalon_anti_slave_0_byteenable;                                        // onchip_memory_s1_translator:av_byteenable -> onchip_memory:byteenable
	wire         ext_flash_uas_translator_avalon_anti_slave_0_waitrequest;                                          // ext_flash:uas_waitrequest -> ext_flash_uas_translator:av_waitrequest
	wire   [1:0] ext_flash_uas_translator_avalon_anti_slave_0_burstcount;                                           // ext_flash_uas_translator:av_burstcount -> ext_flash:uas_burstcount
	wire  [15:0] ext_flash_uas_translator_avalon_anti_slave_0_writedata;                                            // ext_flash_uas_translator:av_writedata -> ext_flash:uas_writedata
	wire  [24:0] ext_flash_uas_translator_avalon_anti_slave_0_address;                                              // ext_flash_uas_translator:av_address -> ext_flash:uas_address
	wire         ext_flash_uas_translator_avalon_anti_slave_0_lock;                                                 // ext_flash_uas_translator:av_lock -> ext_flash:uas_lock
	wire         ext_flash_uas_translator_avalon_anti_slave_0_write;                                                // ext_flash_uas_translator:av_write -> ext_flash:uas_write
	wire         ext_flash_uas_translator_avalon_anti_slave_0_read;                                                 // ext_flash_uas_translator:av_read -> ext_flash:uas_read
	wire  [15:0] ext_flash_uas_translator_avalon_anti_slave_0_readdata;                                             // ext_flash:uas_readdata -> ext_flash_uas_translator:av_readdata
	wire         ext_flash_uas_translator_avalon_anti_slave_0_debugaccess;                                          // ext_flash_uas_translator:av_debugaccess -> ext_flash:uas_debugaccess
	wire         ext_flash_uas_translator_avalon_anti_slave_0_readdatavalid;                                        // ext_flash:uas_readdatavalid -> ext_flash_uas_translator:av_readdatavalid
	wire   [1:0] ext_flash_uas_translator_avalon_anti_slave_0_byteenable;                                           // ext_flash_uas_translator:av_byteenable -> ext_flash:uas_byteenable
	wire         sysid_control_slave_translator_avalon_anti_slave_0_address;                                        // sysid_control_slave_translator:av_address -> sysid:address
	wire  [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                       // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                            // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                              // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                             // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                  // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                   // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                               // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire  [15:0] high_res_timer_s1_translator_avalon_anti_slave_0_writedata;                                        // high_res_timer_s1_translator:av_writedata -> high_res_timer:writedata
	wire   [2:0] high_res_timer_s1_translator_avalon_anti_slave_0_address;                                          // high_res_timer_s1_translator:av_address -> high_res_timer:address
	wire         high_res_timer_s1_translator_avalon_anti_slave_0_chipselect;                                       // high_res_timer_s1_translator:av_chipselect -> high_res_timer:chipselect
	wire         high_res_timer_s1_translator_avalon_anti_slave_0_write;                                            // high_res_timer_s1_translator:av_write -> high_res_timer:write_n
	wire  [15:0] high_res_timer_s1_translator_avalon_anti_slave_0_readdata;                                         // high_res_timer:readdata -> high_res_timer_s1_translator:av_readdata
	wire  [15:0] sys_timer_s1_translator_avalon_anti_slave_0_writedata;                                             // sys_timer_s1_translator:av_writedata -> sys_timer:writedata
	wire   [2:0] sys_timer_s1_translator_avalon_anti_slave_0_address;                                               // sys_timer_s1_translator:av_address -> sys_timer:address
	wire         sys_timer_s1_translator_avalon_anti_slave_0_chipselect;                                            // sys_timer_s1_translator:av_chipselect -> sys_timer:chipselect
	wire         sys_timer_s1_translator_avalon_anti_slave_0_write;                                                 // sys_timer_s1_translator:av_write -> sys_timer:write_n
	wire  [15:0] sys_timer_s1_translator_avalon_anti_slave_0_readdata;                                              // sys_timer:readdata -> sys_timer_s1_translator:av_readdata
	wire         tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest;                                   // tse_mac:waitrequest -> tse_mac_control_port_translator:av_waitrequest
	wire  [31:0] tse_mac_control_port_translator_avalon_anti_slave_0_writedata;                                     // tse_mac_control_port_translator:av_writedata -> tse_mac:writedata
	wire   [7:0] tse_mac_control_port_translator_avalon_anti_slave_0_address;                                       // tse_mac_control_port_translator:av_address -> tse_mac:address
	wire         tse_mac_control_port_translator_avalon_anti_slave_0_write;                                         // tse_mac_control_port_translator:av_write -> tse_mac:write
	wire         tse_mac_control_port_translator_avalon_anti_slave_0_read;                                          // tse_mac_control_port_translator:av_read -> tse_mac:read
	wire  [31:0] tse_mac_control_port_translator_avalon_anti_slave_0_readdata;                                      // tse_mac:readdata -> tse_mac_control_port_translator:av_readdata
	wire  [31:0] sgdma_tx_csr_translator_avalon_anti_slave_0_writedata;                                             // sgdma_tx_csr_translator:av_writedata -> sgdma_tx:csr_writedata
	wire   [3:0] sgdma_tx_csr_translator_avalon_anti_slave_0_address;                                               // sgdma_tx_csr_translator:av_address -> sgdma_tx:csr_address
	wire         sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect;                                            // sgdma_tx_csr_translator:av_chipselect -> sgdma_tx:csr_chipselect
	wire         sgdma_tx_csr_translator_avalon_anti_slave_0_write;                                                 // sgdma_tx_csr_translator:av_write -> sgdma_tx:csr_write
	wire         sgdma_tx_csr_translator_avalon_anti_slave_0_read;                                                  // sgdma_tx_csr_translator:av_read -> sgdma_tx:csr_read
	wire  [31:0] sgdma_tx_csr_translator_avalon_anti_slave_0_readdata;                                              // sgdma_tx:csr_readdata -> sgdma_tx_csr_translator:av_readdata
	wire  [31:0] sgdma_rx_csr_translator_avalon_anti_slave_0_writedata;                                             // sgdma_rx_csr_translator:av_writedata -> sgdma_rx:csr_writedata
	wire   [3:0] sgdma_rx_csr_translator_avalon_anti_slave_0_address;                                               // sgdma_rx_csr_translator:av_address -> sgdma_rx:csr_address
	wire         sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect;                                            // sgdma_rx_csr_translator:av_chipselect -> sgdma_rx:csr_chipselect
	wire         sgdma_rx_csr_translator_avalon_anti_slave_0_write;                                                 // sgdma_rx_csr_translator:av_write -> sgdma_rx:csr_write
	wire         sgdma_rx_csr_translator_avalon_anti_slave_0_read;                                                  // sgdma_rx_csr_translator:av_read -> sgdma_rx:csr_read
	wire  [31:0] sgdma_rx_csr_translator_avalon_anti_slave_0_readdata;                                              // sgdma_rx:csr_readdata -> sgdma_rx_csr_translator:av_readdata
	wire  [31:0] descriptor_memory_s1_translator_avalon_anti_slave_0_writedata;                                     // descriptor_memory_s1_translator:av_writedata -> descriptor_memory:writedata
	wire   [8:0] descriptor_memory_s1_translator_avalon_anti_slave_0_address;                                       // descriptor_memory_s1_translator:av_address -> descriptor_memory:address
	wire         descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect;                                    // descriptor_memory_s1_translator:av_chipselect -> descriptor_memory:chipselect
	wire         descriptor_memory_s1_translator_avalon_anti_slave_0_clken;                                         // descriptor_memory_s1_translator:av_clken -> descriptor_memory:clken
	wire         descriptor_memory_s1_translator_avalon_anti_slave_0_write;                                         // descriptor_memory_s1_translator:av_write -> descriptor_memory:write
	wire  [31:0] descriptor_memory_s1_translator_avalon_anti_slave_0_readdata;                                      // descriptor_memory:readdata -> descriptor_memory_s1_translator:av_readdata
	wire   [3:0] descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable;                                    // descriptor_memory_s1_translator:av_byteenable -> descriptor_memory:byteenable
	wire         peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_waitrequest;                           // peripheral_clock_crossing:s0_waitrequest -> peripheral_clock_crossing_s0_translator:av_waitrequest
	wire         peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_burstcount;                            // peripheral_clock_crossing_s0_translator:av_burstcount -> peripheral_clock_crossing:s0_burstcount
	wire  [31:0] peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_writedata;                             // peripheral_clock_crossing_s0_translator:av_writedata -> peripheral_clock_crossing:s0_writedata
	wire   [5:0] peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_address;                               // peripheral_clock_crossing_s0_translator:av_address -> peripheral_clock_crossing:s0_address
	wire         peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_write;                                 // peripheral_clock_crossing_s0_translator:av_write -> peripheral_clock_crossing:s0_write
	wire         peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_read;                                  // peripheral_clock_crossing_s0_translator:av_read -> peripheral_clock_crossing:s0_read
	wire  [31:0] peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_readdata;                              // peripheral_clock_crossing:s0_readdata -> peripheral_clock_crossing_s0_translator:av_readdata
	wire         peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_debugaccess;                           // peripheral_clock_crossing_s0_translator:av_debugaccess -> peripheral_clock_crossing:s0_debugaccess
	wire         peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_readdatavalid;                         // peripheral_clock_crossing:s0_readdatavalid -> peripheral_clock_crossing_s0_translator:av_readdatavalid
	wire   [3:0] peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_byteenable;                            // peripheral_clock_crossing_s0_translator:av_byteenable -> peripheral_clock_crossing:s0_byteenable
	wire  [31:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata;                                       // altpll_0_pll_slave_translator:av_writedata -> altpll_0:writedata
	wire   [1:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_address;                                         // altpll_0_pll_slave_translator:av_address -> altpll_0:address
	wire         altpll_0_pll_slave_translator_avalon_anti_slave_0_write;                                           // altpll_0_pll_slave_translator:av_write -> altpll_0:write
	wire         altpll_0_pll_slave_translator_avalon_anti_slave_0_read;                                            // altpll_0_pll_slave_translator:av_read -> altpll_0:read
	wire  [31:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata;                                        // altpll_0:readdata -> altpll_0_pll_slave_translator:av_readdata
	wire   [0:0] peripheral_clock_crossing_m0_burstcount;                                                           // peripheral_clock_crossing:m0_burstcount -> peripheral_clock_crossing_m0_translator:av_burstcount
	wire         peripheral_clock_crossing_m0_waitrequest;                                                          // peripheral_clock_crossing_m0_translator:av_waitrequest -> peripheral_clock_crossing:m0_waitrequest
	wire   [5:0] peripheral_clock_crossing_m0_address;                                                              // peripheral_clock_crossing:m0_address -> peripheral_clock_crossing_m0_translator:av_address
	wire  [31:0] peripheral_clock_crossing_m0_writedata;                                                            // peripheral_clock_crossing:m0_writedata -> peripheral_clock_crossing_m0_translator:av_writedata
	wire         peripheral_clock_crossing_m0_write;                                                                // peripheral_clock_crossing:m0_write -> peripheral_clock_crossing_m0_translator:av_write
	wire         peripheral_clock_crossing_m0_read;                                                                 // peripheral_clock_crossing:m0_read -> peripheral_clock_crossing_m0_translator:av_read
	wire  [31:0] peripheral_clock_crossing_m0_readdata;                                                             // peripheral_clock_crossing_m0_translator:av_readdata -> peripheral_clock_crossing:m0_readdata
	wire         peripheral_clock_crossing_m0_debugaccess;                                                          // peripheral_clock_crossing:m0_debugaccess -> peripheral_clock_crossing_m0_translator:av_debugaccess
	wire   [3:0] peripheral_clock_crossing_m0_byteenable;                                                           // peripheral_clock_crossing:m0_byteenable -> peripheral_clock_crossing_m0_translator:av_byteenable
	wire         peripheral_clock_crossing_m0_readdatavalid;                                                        // peripheral_clock_crossing_m0_translator:av_readdatavalid -> peripheral_clock_crossing:m0_readdatavalid
	wire  [31:0] led_pio_s1_translator_avalon_anti_slave_0_writedata;                                               // led_pio_s1_translator:av_writedata -> led_pio:writedata
	wire   [1:0] led_pio_s1_translator_avalon_anti_slave_0_address;                                                 // led_pio_s1_translator:av_address -> led_pio:address
	wire         led_pio_s1_translator_avalon_anti_slave_0_chipselect;                                              // led_pio_s1_translator:av_chipselect -> led_pio:chipselect
	wire         led_pio_s1_translator_avalon_anti_slave_0_write;                                                   // led_pio_s1_translator:av_write -> led_pio:write_n
	wire  [31:0] led_pio_s1_translator_avalon_anti_slave_0_readdata;                                                // led_pio:readdata -> led_pio_s1_translator:av_readdata
	wire   [1:0] sw_pio_s1_translator_avalon_anti_slave_0_address;                                                  // sw_pio_s1_translator:av_address -> sw_pio:address
	wire  [31:0] sw_pio_s1_translator_avalon_anti_slave_0_readdata;                                                 // sw_pio:readdata -> sw_pio_s1_translator:av_readdata
	wire   [1:0] pb_pio_s1_translator_avalon_anti_slave_0_address;                                                  // pb_pio_s1_translator:av_address -> pb_pio:address
	wire  [31:0] pb_pio_s1_translator_avalon_anti_slave_0_readdata;                                                 // pb_pio:readdata -> pb_pio_s1_translator:av_readdata
	wire  [31:0] seven_seg_pio_s1_translator_avalon_anti_slave_0_writedata;                                         // seven_seg_pio_s1_translator:av_writedata -> seven_seg_pio:writedata
	wire   [1:0] seven_seg_pio_s1_translator_avalon_anti_slave_0_address;                                           // seven_seg_pio_s1_translator:av_address -> seven_seg_pio:address
	wire         seven_seg_pio_s1_translator_avalon_anti_slave_0_chipselect;                                        // seven_seg_pio_s1_translator:av_chipselect -> seven_seg_pio:chipselect
	wire         seven_seg_pio_s1_translator_avalon_anti_slave_0_write;                                             // seven_seg_pio_s1_translator:av_write -> seven_seg_pio:write_n
	wire  [31:0] seven_seg_pio_s1_translator_avalon_anti_slave_0_readdata;                                          // seven_seg_pio:readdata -> seven_seg_pio_s1_translator:av_readdata
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // high_res_timer_s1_translator:uav_waitrequest -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> high_res_timer_s1_translator:uav_burstcount
	wire  [31:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> high_res_timer_s1_translator:uav_writedata
	wire  [31:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> high_res_timer_s1_translator:uav_address
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> high_res_timer_s1_translator:uav_write
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> high_res_timer_s1_translator:uav_lock
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> high_res_timer_s1_translator:uav_read
	wire  [31:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // high_res_timer_s1_translator:uav_readdata -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // high_res_timer_s1_translator:uav_readdatavalid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> high_res_timer_s1_translator:uav_debugaccess
	wire   [3:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> high_res_timer_s1_translator:uav_byteenable
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [31:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                  // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                   // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                  // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // cpu_jtag_debug_module_translator:uav_waitrequest -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                      // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_jtag_debug_module_translator:uav_writedata
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_jtag_debug_module_translator:uav_address
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_jtag_debug_module_translator:uav_write
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                           // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_jtag_debug_module_translator:uav_lock
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                           // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                       // cpu_jtag_debug_module_translator:uav_readdata -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // cpu_jtag_debug_module_translator:uav_readdatavalid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_jtag_debug_module_translator:uav_byteenable
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // ext_flash_uas_translator:uav_waitrequest -> ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> ext_flash_uas_translator:uav_burstcount
	wire  [15:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                              // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> ext_flash_uas_translator:uav_writedata
	wire  [31:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_address;                                // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_address -> ext_flash_uas_translator:uav_address
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_write;                                  // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_write -> ext_flash_uas_translator:uav_write
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                   // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_lock -> ext_flash_uas_translator:uav_lock
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_read;                                   // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_read -> ext_flash_uas_translator:uav_read
	wire  [15:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                               // ext_flash_uas_translator:uav_readdata -> ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // ext_flash_uas_translator:uav_readdatavalid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ext_flash_uas_translator:uav_debugaccess
	wire   [1:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> ext_flash_uas_translator:uav_byteenable
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [71:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                            // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [71:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [15:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // peripheral_clock_crossing_s0_translator:uav_waitrequest -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;              // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> peripheral_clock_crossing_s0_translator:uav_burstcount
	wire  [31:0] peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_writedata;               // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> peripheral_clock_crossing_s0_translator:uav_writedata
	wire  [31:0] peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_address;                 // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:m0_address -> peripheral_clock_crossing_s0_translator:uav_address
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_write;                   // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:m0_write -> peripheral_clock_crossing_s0_translator:uav_write
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_lock;                    // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:m0_lock -> peripheral_clock_crossing_s0_translator:uav_lock
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_read;                    // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:m0_read -> peripheral_clock_crossing_s0_translator:uav_read
	wire  [31:0] peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                // peripheral_clock_crossing_s0_translator:uav_readdata -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // peripheral_clock_crossing_s0_translator:uav_readdatavalid -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> peripheral_clock_crossing_s0_translator:uav_debugaccess
	wire   [3:0] peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;              // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> peripheral_clock_crossing_s0_translator:uav_byteenable
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;            // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_data;             // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;            // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest;                                 // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_m_write_translator:uav_waitrequest
	wire   [2:0] sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount;                                  // sgdma_rx_m_write_translator:uav_burstcount -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] sgdma_rx_m_write_translator_avalon_universal_master_0_writedata;                                   // sgdma_rx_m_write_translator:uav_writedata -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] sgdma_rx_m_write_translator_avalon_universal_master_0_address;                                     // sgdma_rx_m_write_translator:uav_address -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_address
	wire         sgdma_rx_m_write_translator_avalon_universal_master_0_lock;                                        // sgdma_rx_m_write_translator:uav_lock -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_lock
	wire         sgdma_rx_m_write_translator_avalon_universal_master_0_write;                                       // sgdma_rx_m_write_translator:uav_write -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_write
	wire         sgdma_rx_m_write_translator_avalon_universal_master_0_read;                                        // sgdma_rx_m_write_translator:uav_read -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] sgdma_rx_m_write_translator_avalon_universal_master_0_readdata;                                    // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_m_write_translator:uav_readdata
	wire         sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess;                                 // sgdma_rx_m_write_translator:uav_debugaccess -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable;                                  // sgdma_rx_m_write_translator:uav_byteenable -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire         sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid;                               // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_m_write_translator:uav_readdatavalid
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // sys_timer_s1_translator:uav_waitrequest -> sys_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // sys_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sys_timer_s1_translator:uav_burstcount
	wire  [31:0] sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // sys_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sys_timer_s1_translator:uav_writedata
	wire  [31:0] sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // sys_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> sys_timer_s1_translator:uav_address
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // sys_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> sys_timer_s1_translator:uav_write
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // sys_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sys_timer_s1_translator:uav_lock
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // sys_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> sys_timer_s1_translator:uav_read
	wire  [31:0] sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // sys_timer_s1_translator:uav_readdata -> sys_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // sys_timer_s1_translator:uav_readdatavalid -> sys_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // sys_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sys_timer_s1_translator:uav_debugaccess
	wire   [3:0] sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // sys_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sys_timer_s1_translator:uav_byteenable
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // sys_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // sys_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // sys_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // sys_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sys_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sys_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sys_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sys_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sys_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // sys_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // sys_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [31:0] sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // sys_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sys_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                       // sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sys_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                        // sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sys_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                       // sys_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire         sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest;                        // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_descriptor_write_translator:uav_waitrequest
	wire   [2:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount;                         // sgdma_rx_descriptor_write_translator:uav_burstcount -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata;                          // sgdma_rx_descriptor_write_translator:uav_writedata -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address;                            // sgdma_rx_descriptor_write_translator:uav_address -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	wire         sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock;                               // sgdma_rx_descriptor_write_translator:uav_lock -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	wire         sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write;                              // sgdma_rx_descriptor_write_translator:uav_write -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	wire         sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read;                               // sgdma_rx_descriptor_write_translator:uav_read -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata;                           // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_descriptor_write_translator:uav_readdata
	wire         sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess;                        // sgdma_rx_descriptor_write_translator:uav_debugaccess -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable;                         // sgdma_rx_descriptor_write_translator:uav_byteenable -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire         sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid;                      // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_descriptor_write_translator:uav_readdatavalid
	wire         sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest;                                  // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_m_read_translator:uav_waitrequest
	wire   [2:0] sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount;                                   // sgdma_tx_m_read_translator:uav_burstcount -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] sgdma_tx_m_read_translator_avalon_universal_master_0_writedata;                                    // sgdma_tx_m_read_translator:uav_writedata -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] sgdma_tx_m_read_translator_avalon_universal_master_0_address;                                      // sgdma_tx_m_read_translator:uav_address -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_address
	wire         sgdma_tx_m_read_translator_avalon_universal_master_0_lock;                                         // sgdma_tx_m_read_translator:uav_lock -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_lock
	wire         sgdma_tx_m_read_translator_avalon_universal_master_0_write;                                        // sgdma_tx_m_read_translator:uav_write -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_write
	wire         sgdma_tx_m_read_translator_avalon_universal_master_0_read;                                         // sgdma_tx_m_read_translator:uav_read -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] sgdma_tx_m_read_translator_avalon_universal_master_0_readdata;                                     // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_m_read_translator:uav_readdata
	wire         sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess;                                  // sgdma_tx_m_read_translator:uav_debugaccess -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable;                                   // sgdma_tx_m_read_translator:uav_byteenable -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire         sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid;                                // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_m_read_translator:uav_readdatavalid
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // sgdma_tx_csr_translator:uav_waitrequest -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> sgdma_tx_csr_translator:uav_burstcount
	wire  [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> sgdma_tx_csr_translator:uav_writedata
	wire  [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_address -> sgdma_tx_csr_translator:uav_address
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_write -> sgdma_tx_csr_translator:uav_write
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_lock -> sgdma_tx_csr_translator:uav_lock
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_read -> sgdma_tx_csr_translator:uav_read
	wire  [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // sgdma_tx_csr_translator:uav_readdata -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // sgdma_tx_csr_translator:uav_readdatavalid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sgdma_tx_csr_translator:uav_debugaccess
	wire   [3:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> sgdma_tx_csr_translator:uav_byteenable
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                         // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire   [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire         sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest;                         // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_descriptor_read_translator:uav_waitrequest
	wire   [2:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount;                          // sgdma_tx_descriptor_read_translator:uav_burstcount -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata;                           // sgdma_tx_descriptor_read_translator:uav_writedata -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address;                             // sgdma_tx_descriptor_read_translator:uav_address -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	wire         sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock;                                // sgdma_tx_descriptor_read_translator:uav_lock -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	wire         sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write;                               // sgdma_tx_descriptor_read_translator:uav_write -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	wire         sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read;                                // sgdma_tx_descriptor_read_translator:uav_read -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata;                            // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_descriptor_read_translator:uav_readdata
	wire         sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess;                         // sgdma_tx_descriptor_read_translator:uav_debugaccess -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable;                          // sgdma_tx_descriptor_read_translator:uav_byteenable -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire         sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid;                       // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_descriptor_read_translator:uav_readdatavalid
	wire         sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest;                        // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_descriptor_write_translator:uav_waitrequest
	wire   [2:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount;                         // sgdma_tx_descriptor_write_translator:uav_burstcount -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata;                          // sgdma_tx_descriptor_write_translator:uav_writedata -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address;                            // sgdma_tx_descriptor_write_translator:uav_address -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	wire         sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock;                               // sgdma_tx_descriptor_write_translator:uav_lock -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	wire         sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write;                              // sgdma_tx_descriptor_write_translator:uav_write -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	wire         sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read;                               // sgdma_tx_descriptor_write_translator:uav_read -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata;                           // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_descriptor_write_translator:uav_readdata
	wire         sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess;                        // sgdma_tx_descriptor_write_translator:uav_debugaccess -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable;                         // sgdma_tx_descriptor_write_translator:uav_byteenable -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire         sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid;                      // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_descriptor_write_translator:uav_readdatavalid
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // tse_mac_control_port_translator:uav_waitrequest -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> tse_mac_control_port_translator:uav_burstcount
	wire  [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;                       // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> tse_mac_control_port_translator:uav_writedata
	wire  [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address;                         // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_address -> tse_mac_control_port_translator:uav_address
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write;                           // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_write -> tse_mac_control_port_translator:uav_write
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                            // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> tse_mac_control_port_translator:uav_lock
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read;                            // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_read -> tse_mac_control_port_translator:uav_read
	wire  [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                        // tse_mac_control_port_translator:uav_readdata -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // tse_mac_control_port_translator:uav_readdatavalid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> tse_mac_control_port_translator:uav_debugaccess
	wire   [3:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> tse_mac_control_port_translator:uav_byteenable
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;                     // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // sgdma_rx_csr_translator:uav_waitrequest -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> sgdma_rx_csr_translator:uav_burstcount
	wire  [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                               // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> sgdma_rx_csr_translator:uav_writedata
	wire  [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address;                                 // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_address -> sgdma_rx_csr_translator:uav_address
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write;                                   // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_write -> sgdma_rx_csr_translator:uav_write
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                    // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_lock -> sgdma_rx_csr_translator:uav_lock
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read;                                    // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_read -> sgdma_rx_csr_translator:uav_read
	wire  [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                // sgdma_rx_csr_translator:uav_readdata -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // sgdma_rx_csr_translator:uav_readdatavalid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sgdma_rx_csr_translator:uav_debugaccess
	wire   [3:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> sgdma_rx_csr_translator:uav_byteenable
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                             // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                           // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                            // cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                             // cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                               // cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_instruction_master_translator_avalon_universal_master_0_lock;                                  // cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_instruction_master_translator_avalon_universal_master_0_write;                                 // cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_instruction_master_translator_avalon_universal_master_0_read;                                  // cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                              // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	wire         cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                           // cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                            // cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                         // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // onchip_memory_s1_translator:uav_waitrequest -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory_s1_translator:uav_burstcount
	wire  [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                           // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory_s1_translator:uav_writedata
	wire  [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                             // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory_s1_translator:uav_address
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                               // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory_s1_translator:uav_write
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory_s1_translator:uav_lock
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                                // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory_s1_translator:uav_read
	wire  [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                            // onchip_memory_s1_translator:uav_readdata -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // onchip_memory_s1_translator:uav_readdatavalid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory_s1_translator:uav_debugaccess
	wire   [3:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory_s1_translator:uav_byteenable
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                         // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // descriptor_memory_s1_translator:uav_waitrequest -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> descriptor_memory_s1_translator:uav_burstcount
	wire  [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                       // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> descriptor_memory_s1_translator:uav_writedata
	wire  [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> descriptor_memory_s1_translator:uav_address
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                           // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> descriptor_memory_s1_translator:uav_write
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                            // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> descriptor_memory_s1_translator:uav_lock
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                            // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> descriptor_memory_s1_translator:uav_read
	wire  [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                        // descriptor_memory_s1_translator:uav_readdata -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // descriptor_memory_s1_translator:uav_readdatavalid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> descriptor_memory_s1_translator:uav_debugaccess
	wire   [3:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> descriptor_memory_s1_translator:uav_byteenable
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                     // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // altpll_0_pll_slave_translator:uav_waitrequest -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> altpll_0_pll_slave_translator:uav_burstcount
	wire  [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                         // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> altpll_0_pll_slave_translator:uav_writedata
	wire  [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                           // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> altpll_0_pll_slave_translator:uav_address
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                             // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> altpll_0_pll_slave_translator:uav_write
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> altpll_0_pll_slave_translator:uav_lock
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> altpll_0_pll_slave_translator:uav_read
	wire  [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                          // altpll_0_pll_slave_translator:uav_readdata -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // altpll_0_pll_slave_translator:uav_readdatavalid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> altpll_0_pll_slave_translator:uav_debugaccess
	wire   [3:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> altpll_0_pll_slave_translator:uav_byteenable
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                       // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                  // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire         sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest;                         // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_descriptor_read_translator:uav_waitrequest
	wire   [2:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount;                          // sgdma_rx_descriptor_read_translator:uav_burstcount -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata;                           // sgdma_rx_descriptor_read_translator:uav_writedata -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address;                             // sgdma_rx_descriptor_read_translator:uav_address -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	wire         sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock;                                // sgdma_rx_descriptor_read_translator:uav_lock -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	wire         sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write;                               // sgdma_rx_descriptor_read_translator:uav_write -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	wire         sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read;                                // sgdma_rx_descriptor_read_translator:uav_read -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata;                            // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_descriptor_read_translator:uav_readdata
	wire         sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess;                         // sgdma_rx_descriptor_read_translator:uav_debugaccess -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable;                          // sgdma_rx_descriptor_read_translator:uav_byteenable -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire         sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid;                       // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_descriptor_read_translator:uav_readdatavalid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                  // cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                   // cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                    // cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] cpu_data_master_translator_avalon_universal_master_0_address;                                      // cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_data_master_translator_avalon_universal_master_0_lock;                                         // cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_data_master_translator_avalon_universal_master_0_write;                                        // cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_data_master_translator_avalon_universal_master_0_read;                                         // cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                     // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	wire         cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                  // cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                   // cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                                // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	wire         peripheral_clock_crossing_m0_translator_avalon_universal_master_0_waitrequest;                     // peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> peripheral_clock_crossing_m0_translator:uav_waitrequest
	wire   [2:0] peripheral_clock_crossing_m0_translator_avalon_universal_master_0_burstcount;                      // peripheral_clock_crossing_m0_translator:uav_burstcount -> peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] peripheral_clock_crossing_m0_translator_avalon_universal_master_0_writedata;                       // peripheral_clock_crossing_m0_translator:uav_writedata -> peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [5:0] peripheral_clock_crossing_m0_translator_avalon_universal_master_0_address;                         // peripheral_clock_crossing_m0_translator:uav_address -> peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:av_address
	wire         peripheral_clock_crossing_m0_translator_avalon_universal_master_0_lock;                            // peripheral_clock_crossing_m0_translator:uav_lock -> peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:av_lock
	wire         peripheral_clock_crossing_m0_translator_avalon_universal_master_0_write;                           // peripheral_clock_crossing_m0_translator:uav_write -> peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:av_write
	wire         peripheral_clock_crossing_m0_translator_avalon_universal_master_0_read;                            // peripheral_clock_crossing_m0_translator:uav_read -> peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] peripheral_clock_crossing_m0_translator_avalon_universal_master_0_readdata;                        // peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:av_readdata -> peripheral_clock_crossing_m0_translator:uav_readdata
	wire         peripheral_clock_crossing_m0_translator_avalon_universal_master_0_debugaccess;                     // peripheral_clock_crossing_m0_translator:uav_debugaccess -> peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] peripheral_clock_crossing_m0_translator_avalon_universal_master_0_byteenable;                      // peripheral_clock_crossing_m0_translator:uav_byteenable -> peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire         peripheral_clock_crossing_m0_translator_avalon_universal_master_0_readdatavalid;                   // peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> peripheral_clock_crossing_m0_translator:uav_readdatavalid
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // seven_seg_pio_s1_translator:uav_waitrequest -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> seven_seg_pio_s1_translator:uav_burstcount
	wire  [31:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                           // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> seven_seg_pio_s1_translator:uav_writedata
	wire   [5:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                             // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> seven_seg_pio_s1_translator:uav_address
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                               // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> seven_seg_pio_s1_translator:uav_write
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> seven_seg_pio_s1_translator:uav_lock
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> seven_seg_pio_s1_translator:uav_read
	wire  [31:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                            // seven_seg_pio_s1_translator:uav_readdata -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // seven_seg_pio_s1_translator:uav_readdatavalid -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> seven_seg_pio_s1_translator:uav_debugaccess
	wire   [3:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> seven_seg_pio_s1_translator:uav_byteenable
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [59:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                         // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [59:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // sw_pio_s1_translator:uav_waitrequest -> sw_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // sw_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sw_pio_s1_translator:uav_burstcount
	wire  [31:0] sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // sw_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sw_pio_s1_translator:uav_writedata
	wire   [5:0] sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // sw_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> sw_pio_s1_translator:uav_address
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // sw_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> sw_pio_s1_translator:uav_write
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // sw_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sw_pio_s1_translator:uav_lock
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // sw_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> sw_pio_s1_translator:uav_read
	wire  [31:0] sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // sw_pio_s1_translator:uav_readdata -> sw_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // sw_pio_s1_translator:uav_readdatavalid -> sw_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // sw_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sw_pio_s1_translator:uav_debugaccess
	wire   [3:0] sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // sw_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sw_pio_s1_translator:uav_byteenable
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // sw_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // sw_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // sw_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [59:0] sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // sw_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sw_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sw_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sw_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sw_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [59:0] sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sw_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // sw_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // sw_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sw_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // sw_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sw_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // sw_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sw_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // led_pio_s1_translator:uav_waitrequest -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_pio_s1_translator:uav_burstcount
	wire  [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_pio_s1_translator:uav_writedata
	wire   [5:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_pio_s1_translator:uav_address
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_pio_s1_translator:uav_write
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_pio_s1_translator:uav_lock
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_pio_s1_translator:uav_read
	wire  [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // led_pio_s1_translator:uav_readdata -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // led_pio_s1_translator:uav_readdatavalid -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_pio_s1_translator:uav_debugaccess
	wire   [3:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_pio_s1_translator:uav_byteenable
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [59:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [59:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // pb_pio_s1_translator:uav_waitrequest -> pb_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // pb_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pb_pio_s1_translator:uav_burstcount
	wire  [31:0] pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // pb_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pb_pio_s1_translator:uav_writedata
	wire   [5:0] pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // pb_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> pb_pio_s1_translator:uav_address
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // pb_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> pb_pio_s1_translator:uav_write
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // pb_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pb_pio_s1_translator:uav_lock
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // pb_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> pb_pio_s1_translator:uav_read
	wire  [31:0] pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // pb_pio_s1_translator:uav_readdata -> pb_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // pb_pio_s1_translator:uav_readdatavalid -> pb_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // pb_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pb_pio_s1_translator:uav_debugaccess
	wire   [3:0] pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // pb_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pb_pio_s1_translator:uav_byteenable
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // pb_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // pb_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // pb_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [59:0] pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // pb_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pb_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pb_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pb_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pb_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [59:0] pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pb_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // pb_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // pb_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pb_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] pb_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // pb_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pb_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // pb_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pb_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                        // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [88:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                         // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                         // cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                               // cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                       // cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [88:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                                // cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                               // addr_router_001:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire         sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid;                      // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire         sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket;              // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [88:0] sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data;                       // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire         sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready;                      // addr_router_002:sink_ready -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	wire         sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket;               // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire         sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid;                     // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire         sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket;             // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [88:0] sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data;                      // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire         sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready;                     // addr_router_003:sink_ready -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	wire         sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire         sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid;                      // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire         sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket;              // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire  [88:0] sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data;                       // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire         sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready;                      // addr_router_004:sink_ready -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	wire         sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket;               // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire         sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid;                     // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire         sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket;             // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire  [88:0] sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data;                      // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire         sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready;                     // addr_router_005:sink_ready -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	wire         sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_006:sink_endofpacket
	wire         sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid;                              // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_006:sink_valid
	wire         sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_006:sink_startofpacket
	wire  [88:0] sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data;                               // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_006:sink_data
	wire         sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_006:sink_ready -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_ready
	wire         sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                         // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_007:sink_endofpacket
	wire         sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid;                               // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_007:sink_valid
	wire         sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket;                       // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_007:sink_startofpacket
	wire  [88:0] sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data;                                // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_007:sink_data
	wire         sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready;                               // addr_router_007:sink_ready -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [88:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                           // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router:sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                               // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [88:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                                // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_001:sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                  // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [70:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_data;                                   // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_002:sink_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [88:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_003:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [88:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_004:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [88:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_005:sink_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // sys_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // sys_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // sys_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [88:0] sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // sys_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_006:sink_ready -> sys_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                           // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [88:0] tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data;                            // tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_007:sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [88:0] sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_008:sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                   // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [88:0] sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data;                                    // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_009:sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                           // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [88:0] descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                            // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire         descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_010:sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_valid;                   // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [88:0] peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_data;                    // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire         peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_011:sink_ready -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                             // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [88:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_012:sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;            // peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_008:sink_endofpacket
	wire         peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_valid;                  // peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_008:sink_valid
	wire         peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;          // peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_008:sink_startofpacket
	wire  [58:0] peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_data;                   // peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_008:sink_data
	wire         peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_ready;                  // addr_router_008:sink_ready -> peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [58:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire         led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_013:sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // sw_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // sw_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // sw_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [58:0] sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // sw_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire         sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_014:sink_ready -> sw_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // pb_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // pb_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // pb_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [58:0] pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // pb_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire         pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_015:sink_ready -> pb_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                               // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [58:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire         seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_016:sink_ready -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                       // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                             // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                     // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [88:0] addr_router_src_data;                                                                              // addr_router:src_data -> limiter:cmd_sink_data
	wire  [12:0] addr_router_src_channel;                                                                           // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                             // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                       // limiter:rsp_src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                             // limiter:rsp_src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                     // limiter:rsp_src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [88:0] limiter_rsp_src_data;                                                                              // limiter:rsp_src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [12:0] limiter_rsp_src_channel;                                                                           // limiter:rsp_src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                             // cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         addr_router_001_src_endofpacket;                                                                   // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire         addr_router_001_src_valid;                                                                         // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire         addr_router_001_src_startofpacket;                                                                 // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [88:0] addr_router_001_src_data;                                                                          // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire  [12:0] addr_router_001_src_channel;                                                                       // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire         addr_router_001_src_ready;                                                                         // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire         limiter_001_rsp_src_endofpacket;                                                                   // limiter_001:rsp_src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_001_rsp_src_valid;                                                                         // limiter_001:rsp_src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_001_rsp_src_startofpacket;                                                                 // limiter_001:rsp_src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [88:0] limiter_001_rsp_src_data;                                                                          // limiter_001:rsp_src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [12:0] limiter_001_rsp_src_channel;                                                                       // limiter_001:rsp_src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_001_rsp_src_ready;                                                                         // cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire         addr_router_002_src_endofpacket;                                                                   // addr_router_002:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	wire         addr_router_002_src_valid;                                                                         // addr_router_002:src_valid -> limiter_002:cmd_sink_valid
	wire         addr_router_002_src_startofpacket;                                                                 // addr_router_002:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	wire  [88:0] addr_router_002_src_data;                                                                          // addr_router_002:src_data -> limiter_002:cmd_sink_data
	wire  [12:0] addr_router_002_src_channel;                                                                       // addr_router_002:src_channel -> limiter_002:cmd_sink_channel
	wire         addr_router_002_src_ready;                                                                         // limiter_002:cmd_sink_ready -> addr_router_002:src_ready
	wire         limiter_002_rsp_src_endofpacket;                                                                   // limiter_002:rsp_src_endofpacket -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_002_rsp_src_valid;                                                                         // limiter_002:rsp_src_valid -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_002_rsp_src_startofpacket;                                                                 // limiter_002:rsp_src_startofpacket -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [88:0] limiter_002_rsp_src_data;                                                                          // limiter_002:rsp_src_data -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	wire  [12:0] limiter_002_rsp_src_channel;                                                                       // limiter_002:rsp_src_channel -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_002_rsp_src_ready;                                                                         // sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	wire         addr_router_004_src_endofpacket;                                                                   // addr_router_004:src_endofpacket -> limiter_003:cmd_sink_endofpacket
	wire         addr_router_004_src_valid;                                                                         // addr_router_004:src_valid -> limiter_003:cmd_sink_valid
	wire         addr_router_004_src_startofpacket;                                                                 // addr_router_004:src_startofpacket -> limiter_003:cmd_sink_startofpacket
	wire  [88:0] addr_router_004_src_data;                                                                          // addr_router_004:src_data -> limiter_003:cmd_sink_data
	wire  [12:0] addr_router_004_src_channel;                                                                       // addr_router_004:src_channel -> limiter_003:cmd_sink_channel
	wire         addr_router_004_src_ready;                                                                         // limiter_003:cmd_sink_ready -> addr_router_004:src_ready
	wire         limiter_003_rsp_src_endofpacket;                                                                   // limiter_003:rsp_src_endofpacket -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_003_rsp_src_valid;                                                                         // limiter_003:rsp_src_valid -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_003_rsp_src_startofpacket;                                                                 // limiter_003:rsp_src_startofpacket -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [88:0] limiter_003_rsp_src_data;                                                                          // limiter_003:rsp_src_data -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	wire  [12:0] limiter_003_rsp_src_channel;                                                                       // limiter_003:rsp_src_channel -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_003_rsp_src_ready;                                                                         // sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> limiter_003:rsp_src_ready
	wire         addr_router_007_src_endofpacket;                                                                   // addr_router_007:src_endofpacket -> limiter_004:cmd_sink_endofpacket
	wire         addr_router_007_src_valid;                                                                         // addr_router_007:src_valid -> limiter_004:cmd_sink_valid
	wire         addr_router_007_src_startofpacket;                                                                 // addr_router_007:src_startofpacket -> limiter_004:cmd_sink_startofpacket
	wire  [88:0] addr_router_007_src_data;                                                                          // addr_router_007:src_data -> limiter_004:cmd_sink_data
	wire  [12:0] addr_router_007_src_channel;                                                                       // addr_router_007:src_channel -> limiter_004:cmd_sink_channel
	wire         addr_router_007_src_ready;                                                                         // limiter_004:cmd_sink_ready -> addr_router_007:src_ready
	wire         limiter_004_rsp_src_endofpacket;                                                                   // limiter_004:rsp_src_endofpacket -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_004_rsp_src_valid;                                                                         // limiter_004:rsp_src_valid -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_004_rsp_src_startofpacket;                                                                 // limiter_004:rsp_src_startofpacket -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [88:0] limiter_004_rsp_src_data;                                                                          // limiter_004:rsp_src_data -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_data
	wire  [12:0] limiter_004_rsp_src_channel;                                                                       // limiter_004:rsp_src_channel -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_004_rsp_src_ready;                                                                         // sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_ready -> limiter_004:rsp_src_ready
	wire         addr_router_008_src_endofpacket;                                                                   // addr_router_008:src_endofpacket -> limiter_005:cmd_sink_endofpacket
	wire         addr_router_008_src_valid;                                                                         // addr_router_008:src_valid -> limiter_005:cmd_sink_valid
	wire         addr_router_008_src_startofpacket;                                                                 // addr_router_008:src_startofpacket -> limiter_005:cmd_sink_startofpacket
	wire  [58:0] addr_router_008_src_data;                                                                          // addr_router_008:src_data -> limiter_005:cmd_sink_data
	wire   [3:0] addr_router_008_src_channel;                                                                       // addr_router_008:src_channel -> limiter_005:cmd_sink_channel
	wire         addr_router_008_src_ready;                                                                         // limiter_005:cmd_sink_ready -> addr_router_008:src_ready
	wire         limiter_005_rsp_src_endofpacket;                                                                   // limiter_005:rsp_src_endofpacket -> peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_005_rsp_src_valid;                                                                         // limiter_005:rsp_src_valid -> peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_005_rsp_src_startofpacket;                                                                 // limiter_005:rsp_src_startofpacket -> peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [58:0] limiter_005_rsp_src_data;                                                                          // limiter_005:rsp_src_data -> peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:rp_data
	wire   [3:0] limiter_005_rsp_src_channel;                                                                       // limiter_005:rsp_src_channel -> peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_005_rsp_src_ready;                                                                         // peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_005:rsp_src_ready
	wire         burst_adapter_source0_endofpacket;                                                                 // burst_adapter:source0_endofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_source0_valid;                                                                       // burst_adapter:source0_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_source0_startofpacket;                                                               // burst_adapter:source0_startofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [70:0] burst_adapter_source0_data;                                                                        // burst_adapter:source0_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_source0_ready;                                                                       // ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire  [12:0] burst_adapter_source0_channel;                                                                     // burst_adapter:source0_channel -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rst_controller_reset_out_reset;                                                                    // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, addr_router_005:reset, addr_router_006:reset, addr_router_007:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_demux_005:reset, cmd_xbar_demux_006:reset, cmd_xbar_demux_007:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_010:reset, cpu:reset_n, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_jtag_debug_module_translator:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:in_reset, crosser_003:in_reset, crosser_004:out_reset, crosser_005:out_reset, crosser_006:out_reset, crosser_007:out_reset, descriptor_memory:reset, descriptor_memory_s1_translator:reset, descriptor_memory_s1_translator_avalon_universal_slave_0_agent:reset, descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ext_flash:reset_reset, ext_flash_uas_translator:reset, ext_flash_uas_translator_avalon_universal_slave_0_agent:reset, ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, flash_tristate_bridge_bridge_0:reset, flash_tristate_bridge_pinSharer_0:reset_reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_004:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, limiter_002:reset, limiter_003:reset, limiter_004:reset, onchip_memory:reset, onchip_memory_s1_translator:reset, onchip_memory_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, peripheral_clock_crossing:s0_reset, peripheral_clock_crossing_s0_translator:reset, peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:reset, peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sgdma_rx:system_reset_n, sgdma_rx_csr_translator:reset, sgdma_rx_csr_translator_avalon_universal_slave_0_agent:reset, sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_rx_descriptor_read_translator:reset, sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:reset, sgdma_rx_descriptor_write_translator:reset, sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:reset, sgdma_rx_m_write_translator:reset, sgdma_rx_m_write_translator_avalon_universal_master_0_agent:reset, sgdma_tx:system_reset_n, sgdma_tx_csr_translator:reset, sgdma_tx_csr_translator_avalon_universal_slave_0_agent:reset, sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_tx_descriptor_read_translator:reset, sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:reset, sgdma_tx_descriptor_write_translator:reset, sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:reset, sgdma_tx_m_read_translator:reset, sgdma_tx_m_read_translator_avalon_universal_master_0_agent:reset, tse_mac:reset, tse_mac_control_port_translator:reset, tse_mac_control_port_translator_avalon_universal_slave_0_agent:reset, tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset]
	wire         cpu_jtag_debug_module_reset_reset;                                                                 // cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                                                // rst_controller_001:reset_out -> [addr_router_008:reset, cmd_xbar_demux_008:reset, crosser:out_reset, crosser_001:out_reset, crosser_002:out_reset, crosser_004:in_reset, crosser_005:in_reset, crosser_006:in_reset, high_res_timer:reset_n, high_res_timer_s1_translator:reset, high_res_timer_s1_translator_avalon_universal_slave_0_agent:reset, high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_003:reset, id_router_005:reset, id_router_006:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, led_pio:reset_n, led_pio_s1_translator:reset, led_pio_s1_translator_avalon_universal_slave_0_agent:reset, led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter_005:reset, pb_pio:reset_n, pb_pio_s1_translator:reset, pb_pio_s1_translator_avalon_universal_slave_0_agent:reset, pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, peripheral_clock_crossing:m0_reset, peripheral_clock_crossing_m0_translator:reset, peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_mux_008:reset, seven_seg_pio:reset_n, seven_seg_pio_s1_translator:reset, seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:reset, seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sw_pio:reset_n, sw_pio_s1_translator:reset, sw_pio_s1_translator_avalon_universal_slave_0_agent:reset, sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sys_timer:reset_n, sys_timer_s1_translator:reset, sys_timer_s1_translator_avalon_universal_slave_0_agent:reset, sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         rst_controller_002_reset_out_reset;                                                                // rst_controller_002:reset_out -> [altpll_0:reset, altpll_0_pll_slave_translator:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser_003:out_reset, crosser_007:in_reset, id_router_012:reset, rsp_xbar_demux_012:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                                   // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                         // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                 // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [88:0] cmd_xbar_demux_src0_data;                                                                          // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire  [12:0] cmd_xbar_demux_src0_channel;                                                                       // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                         // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                   // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                         // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                 // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [88:0] cmd_xbar_demux_src1_data;                                                                          // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire  [12:0] cmd_xbar_demux_src1_channel;                                                                       // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                         // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                   // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                         // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                 // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [88:0] cmd_xbar_demux_src2_data;                                                                          // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire  [12:0] cmd_xbar_demux_src2_channel;                                                                       // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                         // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                               // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                     // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                             // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src0_data;                                                                      // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire  [12:0] cmd_xbar_demux_001_src0_channel;                                                                   // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                     // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                               // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                     // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                             // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src1_data;                                                                      // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire  [12:0] cmd_xbar_demux_001_src1_channel;                                                                   // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                     // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                               // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                     // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                             // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src2_data;                                                                      // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire  [12:0] cmd_xbar_demux_001_src2_channel;                                                                   // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                     // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                               // cmd_xbar_demux_001:src4_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                     // cmd_xbar_demux_001:src4_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                             // cmd_xbar_demux_001:src4_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src4_data;                                                                      // cmd_xbar_demux_001:src4_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_demux_001_src4_channel;                                                                   // cmd_xbar_demux_001:src4_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                               // cmd_xbar_demux_001:src7_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                     // cmd_xbar_demux_001:src7_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                             // cmd_xbar_demux_001:src7_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src7_data;                                                                      // cmd_xbar_demux_001:src7_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_demux_001_src7_channel;                                                                   // cmd_xbar_demux_001:src7_channel -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                               // cmd_xbar_demux_001:src8_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                     // cmd_xbar_demux_001:src8_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                             // cmd_xbar_demux_001:src8_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src8_data;                                                                      // cmd_xbar_demux_001:src8_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_demux_001_src8_channel;                                                                   // cmd_xbar_demux_001:src8_channel -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src9_endofpacket;                                                               // cmd_xbar_demux_001:src9_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src9_valid;                                                                     // cmd_xbar_demux_001:src9_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src9_startofpacket;                                                             // cmd_xbar_demux_001:src9_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src9_data;                                                                      // cmd_xbar_demux_001:src9_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_demux_001_src9_channel;                                                                   // cmd_xbar_demux_001:src9_channel -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src10_endofpacket;                                                              // cmd_xbar_demux_001:src10_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	wire         cmd_xbar_demux_001_src10_valid;                                                                    // cmd_xbar_demux_001:src10_valid -> cmd_xbar_mux_010:sink0_valid
	wire         cmd_xbar_demux_001_src10_startofpacket;                                                            // cmd_xbar_demux_001:src10_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src10_data;                                                                     // cmd_xbar_demux_001:src10_data -> cmd_xbar_mux_010:sink0_data
	wire  [12:0] cmd_xbar_demux_001_src10_channel;                                                                  // cmd_xbar_demux_001:src10_channel -> cmd_xbar_mux_010:sink0_channel
	wire         cmd_xbar_demux_001_src10_ready;                                                                    // cmd_xbar_mux_010:sink0_ready -> cmd_xbar_demux_001:src10_ready
	wire         cmd_xbar_demux_001_src11_endofpacket;                                                              // cmd_xbar_demux_001:src11_endofpacket -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src11_valid;                                                                    // cmd_xbar_demux_001:src11_valid -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src11_startofpacket;                                                            // cmd_xbar_demux_001:src11_startofpacket -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src11_data;                                                                     // cmd_xbar_demux_001:src11_data -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_demux_001_src11_channel;                                                                  // cmd_xbar_demux_001:src11_channel -> peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src0_endofpacket;                                                               // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	wire         cmd_xbar_demux_002_src0_valid;                                                                     // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_010:sink1_valid
	wire         cmd_xbar_demux_002_src0_startofpacket;                                                             // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	wire  [88:0] cmd_xbar_demux_002_src0_data;                                                                      // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_010:sink1_data
	wire  [12:0] cmd_xbar_demux_002_src0_channel;                                                                   // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_010:sink1_channel
	wire         cmd_xbar_demux_002_src0_ready;                                                                     // cmd_xbar_mux_010:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire         cmd_xbar_demux_003_src0_endofpacket;                                                               // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_010:sink2_endofpacket
	wire         cmd_xbar_demux_003_src0_valid;                                                                     // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_010:sink2_valid
	wire         cmd_xbar_demux_003_src0_startofpacket;                                                             // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_010:sink2_startofpacket
	wire  [88:0] cmd_xbar_demux_003_src0_data;                                                                      // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_010:sink2_data
	wire  [12:0] cmd_xbar_demux_003_src0_channel;                                                                   // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_010:sink2_channel
	wire         cmd_xbar_demux_003_src0_ready;                                                                     // cmd_xbar_mux_010:sink2_ready -> cmd_xbar_demux_003:src0_ready
	wire         cmd_xbar_demux_004_src0_endofpacket;                                                               // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_010:sink3_endofpacket
	wire         cmd_xbar_demux_004_src0_valid;                                                                     // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_010:sink3_valid
	wire         cmd_xbar_demux_004_src0_startofpacket;                                                             // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_010:sink3_startofpacket
	wire  [88:0] cmd_xbar_demux_004_src0_data;                                                                      // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_010:sink3_data
	wire  [12:0] cmd_xbar_demux_004_src0_channel;                                                                   // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_010:sink3_channel
	wire         cmd_xbar_demux_004_src0_ready;                                                                     // cmd_xbar_mux_010:sink3_ready -> cmd_xbar_demux_004:src0_ready
	wire         cmd_xbar_demux_005_src0_endofpacket;                                                               // cmd_xbar_demux_005:src0_endofpacket -> cmd_xbar_mux_010:sink4_endofpacket
	wire         cmd_xbar_demux_005_src0_valid;                                                                     // cmd_xbar_demux_005:src0_valid -> cmd_xbar_mux_010:sink4_valid
	wire         cmd_xbar_demux_005_src0_startofpacket;                                                             // cmd_xbar_demux_005:src0_startofpacket -> cmd_xbar_mux_010:sink4_startofpacket
	wire  [88:0] cmd_xbar_demux_005_src0_data;                                                                      // cmd_xbar_demux_005:src0_data -> cmd_xbar_mux_010:sink4_data
	wire  [12:0] cmd_xbar_demux_005_src0_channel;                                                                   // cmd_xbar_demux_005:src0_channel -> cmd_xbar_mux_010:sink4_channel
	wire         cmd_xbar_demux_005_src0_ready;                                                                     // cmd_xbar_mux_010:sink4_ready -> cmd_xbar_demux_005:src0_ready
	wire         cmd_xbar_demux_006_src0_endofpacket;                                                               // cmd_xbar_demux_006:src0_endofpacket -> cmd_xbar_mux_001:sink2_endofpacket
	wire         cmd_xbar_demux_006_src0_valid;                                                                     // cmd_xbar_demux_006:src0_valid -> cmd_xbar_mux_001:sink2_valid
	wire         cmd_xbar_demux_006_src0_startofpacket;                                                             // cmd_xbar_demux_006:src0_startofpacket -> cmd_xbar_mux_001:sink2_startofpacket
	wire  [88:0] cmd_xbar_demux_006_src0_data;                                                                      // cmd_xbar_demux_006:src0_data -> cmd_xbar_mux_001:sink2_data
	wire  [12:0] cmd_xbar_demux_006_src0_channel;                                                                   // cmd_xbar_demux_006:src0_channel -> cmd_xbar_mux_001:sink2_channel
	wire         cmd_xbar_demux_006_src0_ready;                                                                     // cmd_xbar_mux_001:sink2_ready -> cmd_xbar_demux_006:src0_ready
	wire         cmd_xbar_demux_007_src0_endofpacket;                                                               // cmd_xbar_demux_007:src0_endofpacket -> cmd_xbar_mux_001:sink3_endofpacket
	wire         cmd_xbar_demux_007_src0_valid;                                                                     // cmd_xbar_demux_007:src0_valid -> cmd_xbar_mux_001:sink3_valid
	wire         cmd_xbar_demux_007_src0_startofpacket;                                                             // cmd_xbar_demux_007:src0_startofpacket -> cmd_xbar_mux_001:sink3_startofpacket
	wire  [88:0] cmd_xbar_demux_007_src0_data;                                                                      // cmd_xbar_demux_007:src0_data -> cmd_xbar_mux_001:sink3_data
	wire  [12:0] cmd_xbar_demux_007_src0_channel;                                                                   // cmd_xbar_demux_007:src0_channel -> cmd_xbar_mux_001:sink3_channel
	wire         cmd_xbar_demux_007_src0_ready;                                                                     // cmd_xbar_mux_001:sink3_ready -> cmd_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_src0_endofpacket;                                                                   // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                         // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                 // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [88:0] rsp_xbar_demux_src0_data;                                                                          // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire  [12:0] rsp_xbar_demux_src0_channel;                                                                       // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                         // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                   // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                         // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                 // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [88:0] rsp_xbar_demux_src1_data;                                                                          // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire  [12:0] rsp_xbar_demux_src1_channel;                                                                       // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                         // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                               // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                     // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                             // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [88:0] rsp_xbar_demux_001_src0_data;                                                                      // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire  [12:0] rsp_xbar_demux_001_src0_channel;                                                                   // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                     // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                               // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                     // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                             // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [88:0] rsp_xbar_demux_001_src1_data;                                                                      // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire  [12:0] rsp_xbar_demux_001_src1_channel;                                                                   // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                     // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_001_src2_endofpacket;                                                               // rsp_xbar_demux_001:src2_endofpacket -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_001_src2_valid;                                                                     // rsp_xbar_demux_001:src2_valid -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_001_src2_startofpacket;                                                             // rsp_xbar_demux_001:src2_startofpacket -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [88:0] rsp_xbar_demux_001_src2_data;                                                                      // rsp_xbar_demux_001:src2_data -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_data
	wire  [12:0] rsp_xbar_demux_001_src2_channel;                                                                   // rsp_xbar_demux_001:src2_channel -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_demux_001_src3_endofpacket;                                                               // rsp_xbar_demux_001:src3_endofpacket -> limiter_004:rsp_sink_endofpacket
	wire         rsp_xbar_demux_001_src3_valid;                                                                     // rsp_xbar_demux_001:src3_valid -> limiter_004:rsp_sink_valid
	wire         rsp_xbar_demux_001_src3_startofpacket;                                                             // rsp_xbar_demux_001:src3_startofpacket -> limiter_004:rsp_sink_startofpacket
	wire  [88:0] rsp_xbar_demux_001_src3_data;                                                                      // rsp_xbar_demux_001:src3_data -> limiter_004:rsp_sink_data
	wire  [12:0] rsp_xbar_demux_001_src3_channel;                                                                   // rsp_xbar_demux_001:src3_channel -> limiter_004:rsp_sink_channel
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                               // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                     // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                             // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [88:0] rsp_xbar_demux_002_src0_data;                                                                      // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire  [12:0] rsp_xbar_demux_002_src0_channel;                                                                   // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                     // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                               // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                     // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                             // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [88:0] rsp_xbar_demux_002_src1_data;                                                                      // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire  [12:0] rsp_xbar_demux_002_src1_channel;                                                                   // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                     // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                               // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                     // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                             // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [88:0] rsp_xbar_demux_004_src0_data;                                                                      // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire  [12:0] rsp_xbar_demux_004_src0_channel;                                                                   // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                     // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                               // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                     // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                             // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [88:0] rsp_xbar_demux_007_src0_data;                                                                      // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire  [12:0] rsp_xbar_demux_007_src0_channel;                                                                   // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                     // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                               // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                     // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                             // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [88:0] rsp_xbar_demux_008_src0_data;                                                                      // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire  [12:0] rsp_xbar_demux_008_src0_channel;                                                                   // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                     // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                               // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                                     // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                             // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [88:0] rsp_xbar_demux_009_src0_data;                                                                      // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire  [12:0] rsp_xbar_demux_009_src0_channel;                                                                   // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                                     // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire         rsp_xbar_demux_010_src0_endofpacket;                                                               // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire         rsp_xbar_demux_010_src0_valid;                                                                     // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire         rsp_xbar_demux_010_src0_startofpacket;                                                             // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [88:0] rsp_xbar_demux_010_src0_data;                                                                      // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire  [12:0] rsp_xbar_demux_010_src0_channel;                                                                   // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire         rsp_xbar_demux_010_src0_ready;                                                                     // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire         rsp_xbar_demux_010_src1_endofpacket;                                                               // rsp_xbar_demux_010:src1_endofpacket -> limiter_002:rsp_sink_endofpacket
	wire         rsp_xbar_demux_010_src1_valid;                                                                     // rsp_xbar_demux_010:src1_valid -> limiter_002:rsp_sink_valid
	wire         rsp_xbar_demux_010_src1_startofpacket;                                                             // rsp_xbar_demux_010:src1_startofpacket -> limiter_002:rsp_sink_startofpacket
	wire  [88:0] rsp_xbar_demux_010_src1_data;                                                                      // rsp_xbar_demux_010:src1_data -> limiter_002:rsp_sink_data
	wire  [12:0] rsp_xbar_demux_010_src1_channel;                                                                   // rsp_xbar_demux_010:src1_channel -> limiter_002:rsp_sink_channel
	wire         rsp_xbar_demux_010_src2_endofpacket;                                                               // rsp_xbar_demux_010:src2_endofpacket -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_010_src2_valid;                                                                     // rsp_xbar_demux_010:src2_valid -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_010_src2_startofpacket;                                                             // rsp_xbar_demux_010:src2_startofpacket -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [88:0] rsp_xbar_demux_010_src2_data;                                                                      // rsp_xbar_demux_010:src2_data -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	wire  [12:0] rsp_xbar_demux_010_src2_channel;                                                                   // rsp_xbar_demux_010:src2_channel -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_demux_010_src3_endofpacket;                                                               // rsp_xbar_demux_010:src3_endofpacket -> limiter_003:rsp_sink_endofpacket
	wire         rsp_xbar_demux_010_src3_valid;                                                                     // rsp_xbar_demux_010:src3_valid -> limiter_003:rsp_sink_valid
	wire         rsp_xbar_demux_010_src3_startofpacket;                                                             // rsp_xbar_demux_010:src3_startofpacket -> limiter_003:rsp_sink_startofpacket
	wire  [88:0] rsp_xbar_demux_010_src3_data;                                                                      // rsp_xbar_demux_010:src3_data -> limiter_003:rsp_sink_data
	wire  [12:0] rsp_xbar_demux_010_src3_channel;                                                                   // rsp_xbar_demux_010:src3_channel -> limiter_003:rsp_sink_channel
	wire         rsp_xbar_demux_010_src4_endofpacket;                                                               // rsp_xbar_demux_010:src4_endofpacket -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_010_src4_valid;                                                                     // rsp_xbar_demux_010:src4_valid -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_010_src4_startofpacket;                                                             // rsp_xbar_demux_010:src4_startofpacket -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [88:0] rsp_xbar_demux_010_src4_data;                                                                      // rsp_xbar_demux_010:src4_data -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	wire  [12:0] rsp_xbar_demux_010_src4_channel;                                                                   // rsp_xbar_demux_010:src4_channel -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_demux_011_src0_endofpacket;                                                               // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire         rsp_xbar_demux_011_src0_valid;                                                                     // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire         rsp_xbar_demux_011_src0_startofpacket;                                                             // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [88:0] rsp_xbar_demux_011_src0_data;                                                                      // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire  [12:0] rsp_xbar_demux_011_src0_channel;                                                                   // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire         rsp_xbar_demux_011_src0_ready;                                                                     // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                       // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                     // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [88:0] limiter_cmd_src_data;                                                                              // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire  [12:0] limiter_cmd_src_channel;                                                                           // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                             // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                      // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                            // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                    // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [88:0] rsp_xbar_mux_src_data;                                                                             // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire  [12:0] rsp_xbar_mux_src_channel;                                                                          // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                            // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         limiter_001_cmd_src_endofpacket;                                                                   // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         limiter_001_cmd_src_startofpacket;                                                                 // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [88:0] limiter_001_cmd_src_data;                                                                          // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire  [12:0] limiter_001_cmd_src_channel;                                                                       // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire         limiter_001_cmd_src_ready;                                                                         // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                  // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                        // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [88:0] rsp_xbar_mux_001_src_data;                                                                         // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire  [12:0] rsp_xbar_mux_001_src_channel;                                                                      // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                        // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire         limiter_002_cmd_src_endofpacket;                                                                   // limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire         limiter_002_cmd_src_startofpacket;                                                                 // limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [88:0] limiter_002_cmd_src_data;                                                                          // limiter_002:cmd_src_data -> cmd_xbar_demux_002:sink_data
	wire  [12:0] limiter_002_cmd_src_channel;                                                                       // limiter_002:cmd_src_channel -> cmd_xbar_demux_002:sink_channel
	wire         limiter_002_cmd_src_ready;                                                                         // cmd_xbar_demux_002:sink_ready -> limiter_002:cmd_src_ready
	wire         rsp_xbar_demux_010_src1_ready;                                                                     // limiter_002:rsp_sink_ready -> rsp_xbar_demux_010:src1_ready
	wire         addr_router_003_src_endofpacket;                                                                   // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire         addr_router_003_src_valid;                                                                         // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire         addr_router_003_src_startofpacket;                                                                 // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [88:0] addr_router_003_src_data;                                                                          // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire  [12:0] addr_router_003_src_channel;                                                                       // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire         addr_router_003_src_ready;                                                                         // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire         rsp_xbar_demux_010_src2_ready;                                                                     // sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_010:src2_ready
	wire         limiter_003_cmd_src_endofpacket;                                                                   // limiter_003:cmd_src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire         limiter_003_cmd_src_startofpacket;                                                                 // limiter_003:cmd_src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire  [88:0] limiter_003_cmd_src_data;                                                                          // limiter_003:cmd_src_data -> cmd_xbar_demux_004:sink_data
	wire  [12:0] limiter_003_cmd_src_channel;                                                                       // limiter_003:cmd_src_channel -> cmd_xbar_demux_004:sink_channel
	wire         limiter_003_cmd_src_ready;                                                                         // cmd_xbar_demux_004:sink_ready -> limiter_003:cmd_src_ready
	wire         rsp_xbar_demux_010_src3_ready;                                                                     // limiter_003:rsp_sink_ready -> rsp_xbar_demux_010:src3_ready
	wire         addr_router_005_src_endofpacket;                                                                   // addr_router_005:src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire         addr_router_005_src_valid;                                                                         // addr_router_005:src_valid -> cmd_xbar_demux_005:sink_valid
	wire         addr_router_005_src_startofpacket;                                                                 // addr_router_005:src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire  [88:0] addr_router_005_src_data;                                                                          // addr_router_005:src_data -> cmd_xbar_demux_005:sink_data
	wire  [12:0] addr_router_005_src_channel;                                                                       // addr_router_005:src_channel -> cmd_xbar_demux_005:sink_channel
	wire         addr_router_005_src_ready;                                                                         // cmd_xbar_demux_005:sink_ready -> addr_router_005:src_ready
	wire         rsp_xbar_demux_010_src4_ready;                                                                     // sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_010:src4_ready
	wire         addr_router_006_src_endofpacket;                                                                   // addr_router_006:src_endofpacket -> cmd_xbar_demux_006:sink_endofpacket
	wire         addr_router_006_src_valid;                                                                         // addr_router_006:src_valid -> cmd_xbar_demux_006:sink_valid
	wire         addr_router_006_src_startofpacket;                                                                 // addr_router_006:src_startofpacket -> cmd_xbar_demux_006:sink_startofpacket
	wire  [88:0] addr_router_006_src_data;                                                                          // addr_router_006:src_data -> cmd_xbar_demux_006:sink_data
	wire  [12:0] addr_router_006_src_channel;                                                                       // addr_router_006:src_channel -> cmd_xbar_demux_006:sink_channel
	wire         addr_router_006_src_ready;                                                                         // cmd_xbar_demux_006:sink_ready -> addr_router_006:src_ready
	wire         rsp_xbar_demux_001_src2_ready;                                                                     // sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_001:src2_ready
	wire         limiter_004_cmd_src_endofpacket;                                                                   // limiter_004:cmd_src_endofpacket -> cmd_xbar_demux_007:sink_endofpacket
	wire         limiter_004_cmd_src_startofpacket;                                                                 // limiter_004:cmd_src_startofpacket -> cmd_xbar_demux_007:sink_startofpacket
	wire  [88:0] limiter_004_cmd_src_data;                                                                          // limiter_004:cmd_src_data -> cmd_xbar_demux_007:sink_data
	wire  [12:0] limiter_004_cmd_src_channel;                                                                       // limiter_004:cmd_src_channel -> cmd_xbar_demux_007:sink_channel
	wire         limiter_004_cmd_src_ready;                                                                         // cmd_xbar_demux_007:sink_ready -> limiter_004:cmd_src_ready
	wire         rsp_xbar_demux_001_src3_ready;                                                                     // limiter_004:rsp_sink_ready -> rsp_xbar_demux_001:src3_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                      // cmd_xbar_mux:src_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                            // cmd_xbar_mux:src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                    // cmd_xbar_mux:src_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] cmd_xbar_mux_src_data;                                                                             // cmd_xbar_mux:src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_mux_src_channel;                                                                          // cmd_xbar_mux:src_channel -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                         // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                               // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                       // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [88:0] id_router_src_data;                                                                                // id_router:src_data -> rsp_xbar_demux:sink_data
	wire  [12:0] id_router_src_channel;                                                                             // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                               // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                  // cmd_xbar_mux_001:src_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                        // cmd_xbar_mux_001:src_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                // cmd_xbar_mux_001:src_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] cmd_xbar_mux_001_src_data;                                                                         // cmd_xbar_mux_001:src_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_mux_001_src_channel;                                                                      // cmd_xbar_mux_001:src_channel -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                        // onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                     // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                           // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                   // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [88:0] id_router_001_src_data;                                                                            // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire  [12:0] id_router_001_src_channel;                                                                         // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                           // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         crosser_out_ready;                                                                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire         id_router_003_src_endofpacket;                                                                     // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                           // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                   // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [88:0] id_router_003_src_data;                                                                            // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire  [12:0] id_router_003_src_channel;                                                                         // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                           // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_001_src4_ready;                                                                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire         id_router_004_src_endofpacket;                                                                     // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                           // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                   // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [88:0] id_router_004_src_data;                                                                            // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire  [12:0] id_router_004_src_channel;                                                                         // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                           // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         crosser_001_out_ready;                                                                             // high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_001:out_ready
	wire         id_router_005_src_endofpacket;                                                                     // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                           // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                   // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [88:0] id_router_005_src_data;                                                                            // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire  [12:0] id_router_005_src_channel;                                                                         // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                           // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         crosser_002_out_ready;                                                                             // sys_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_002:out_ready
	wire         id_router_006_src_endofpacket;                                                                     // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                           // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                   // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [88:0] id_router_006_src_data;                                                                            // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire  [12:0] id_router_006_src_channel;                                                                         // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                           // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_demux_001_src7_ready;                                                                     // tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire         id_router_007_src_endofpacket;                                                                     // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                           // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                   // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [88:0] id_router_007_src_data;                                                                            // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire  [12:0] id_router_007_src_channel;                                                                         // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                           // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_demux_001_src8_ready;                                                                     // sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire         id_router_008_src_endofpacket;                                                                     // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                           // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                   // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [88:0] id_router_008_src_data;                                                                            // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire  [12:0] id_router_008_src_channel;                                                                         // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                           // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_demux_001_src9_ready;                                                                     // sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire         id_router_009_src_endofpacket;                                                                     // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         id_router_009_src_valid;                                                                           // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire         id_router_009_src_startofpacket;                                                                   // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [88:0] id_router_009_src_data;                                                                            // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire  [12:0] id_router_009_src_channel;                                                                         // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire         id_router_009_src_ready;                                                                           // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire         cmd_xbar_mux_010_src_endofpacket;                                                                  // cmd_xbar_mux_010:src_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_010_src_valid;                                                                        // cmd_xbar_mux_010:src_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_010_src_startofpacket;                                                                // cmd_xbar_mux_010:src_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] cmd_xbar_mux_010_src_data;                                                                         // cmd_xbar_mux_010:src_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] cmd_xbar_mux_010_src_channel;                                                                      // cmd_xbar_mux_010:src_channel -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_010_src_ready;                                                                        // descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_010:src_ready
	wire         id_router_010_src_endofpacket;                                                                     // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire         id_router_010_src_valid;                                                                           // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire         id_router_010_src_startofpacket;                                                                   // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [88:0] id_router_010_src_data;                                                                            // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire  [12:0] id_router_010_src_channel;                                                                         // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire         id_router_010_src_ready;                                                                           // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire         cmd_xbar_demux_001_src11_ready;                                                                    // peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire         id_router_011_src_endofpacket;                                                                     // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire         id_router_011_src_valid;                                                                           // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire         id_router_011_src_startofpacket;                                                                   // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [88:0] id_router_011_src_data;                                                                            // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire  [12:0] id_router_011_src_channel;                                                                         // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire         id_router_011_src_ready;                                                                           // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire         crosser_003_out_ready;                                                                             // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_003:out_ready
	wire         id_router_012_src_endofpacket;                                                                     // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire         id_router_012_src_valid;                                                                           // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire         id_router_012_src_startofpacket;                                                                   // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [88:0] id_router_012_src_data;                                                                            // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire  [12:0] id_router_012_src_channel;                                                                         // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire         id_router_012_src_ready;                                                                           // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire         cmd_xbar_demux_008_src0_endofpacket;                                                               // cmd_xbar_demux_008:src0_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_008_src0_valid;                                                                     // cmd_xbar_demux_008:src0_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_008_src0_startofpacket;                                                             // cmd_xbar_demux_008:src0_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [58:0] cmd_xbar_demux_008_src0_data;                                                                      // cmd_xbar_demux_008:src0_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [3:0] cmd_xbar_demux_008_src0_channel;                                                                   // cmd_xbar_demux_008:src0_channel -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_008_src1_endofpacket;                                                               // cmd_xbar_demux_008:src1_endofpacket -> sw_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_008_src1_valid;                                                                     // cmd_xbar_demux_008:src1_valid -> sw_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_008_src1_startofpacket;                                                             // cmd_xbar_demux_008:src1_startofpacket -> sw_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [58:0] cmd_xbar_demux_008_src1_data;                                                                      // cmd_xbar_demux_008:src1_data -> sw_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [3:0] cmd_xbar_demux_008_src1_channel;                                                                   // cmd_xbar_demux_008:src1_channel -> sw_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_008_src2_endofpacket;                                                               // cmd_xbar_demux_008:src2_endofpacket -> pb_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_008_src2_valid;                                                                     // cmd_xbar_demux_008:src2_valid -> pb_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_008_src2_startofpacket;                                                             // cmd_xbar_demux_008:src2_startofpacket -> pb_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [58:0] cmd_xbar_demux_008_src2_data;                                                                      // cmd_xbar_demux_008:src2_data -> pb_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [3:0] cmd_xbar_demux_008_src2_channel;                                                                   // cmd_xbar_demux_008:src2_channel -> pb_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_008_src3_endofpacket;                                                               // cmd_xbar_demux_008:src3_endofpacket -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_008_src3_valid;                                                                     // cmd_xbar_demux_008:src3_valid -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_008_src3_startofpacket;                                                             // cmd_xbar_demux_008:src3_startofpacket -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [58:0] cmd_xbar_demux_008_src3_data;                                                                      // cmd_xbar_demux_008:src3_data -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [3:0] cmd_xbar_demux_008_src3_channel;                                                                   // cmd_xbar_demux_008:src3_channel -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_013_src0_endofpacket;                                                               // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_008:sink0_endofpacket
	wire         rsp_xbar_demux_013_src0_valid;                                                                     // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_008:sink0_valid
	wire         rsp_xbar_demux_013_src0_startofpacket;                                                             // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_008:sink0_startofpacket
	wire  [58:0] rsp_xbar_demux_013_src0_data;                                                                      // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_008:sink0_data
	wire   [3:0] rsp_xbar_demux_013_src0_channel;                                                                   // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_008:sink0_channel
	wire         rsp_xbar_demux_013_src0_ready;                                                                     // rsp_xbar_mux_008:sink0_ready -> rsp_xbar_demux_013:src0_ready
	wire         rsp_xbar_demux_014_src0_endofpacket;                                                               // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_008:sink1_endofpacket
	wire         rsp_xbar_demux_014_src0_valid;                                                                     // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_008:sink1_valid
	wire         rsp_xbar_demux_014_src0_startofpacket;                                                             // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_008:sink1_startofpacket
	wire  [58:0] rsp_xbar_demux_014_src0_data;                                                                      // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_008:sink1_data
	wire   [3:0] rsp_xbar_demux_014_src0_channel;                                                                   // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_008:sink1_channel
	wire         rsp_xbar_demux_014_src0_ready;                                                                     // rsp_xbar_mux_008:sink1_ready -> rsp_xbar_demux_014:src0_ready
	wire         rsp_xbar_demux_015_src0_endofpacket;                                                               // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_008:sink2_endofpacket
	wire         rsp_xbar_demux_015_src0_valid;                                                                     // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_008:sink2_valid
	wire         rsp_xbar_demux_015_src0_startofpacket;                                                             // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_008:sink2_startofpacket
	wire  [58:0] rsp_xbar_demux_015_src0_data;                                                                      // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_008:sink2_data
	wire   [3:0] rsp_xbar_demux_015_src0_channel;                                                                   // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_008:sink2_channel
	wire         rsp_xbar_demux_015_src0_ready;                                                                     // rsp_xbar_mux_008:sink2_ready -> rsp_xbar_demux_015:src0_ready
	wire         rsp_xbar_demux_016_src0_endofpacket;                                                               // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_008:sink3_endofpacket
	wire         rsp_xbar_demux_016_src0_valid;                                                                     // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_008:sink3_valid
	wire         rsp_xbar_demux_016_src0_startofpacket;                                                             // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_008:sink3_startofpacket
	wire  [58:0] rsp_xbar_demux_016_src0_data;                                                                      // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_008:sink3_data
	wire   [3:0] rsp_xbar_demux_016_src0_channel;                                                                   // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_008:sink3_channel
	wire         rsp_xbar_demux_016_src0_ready;                                                                     // rsp_xbar_mux_008:sink3_ready -> rsp_xbar_demux_016:src0_ready
	wire         limiter_005_cmd_src_endofpacket;                                                                   // limiter_005:cmd_src_endofpacket -> cmd_xbar_demux_008:sink_endofpacket
	wire         limiter_005_cmd_src_startofpacket;                                                                 // limiter_005:cmd_src_startofpacket -> cmd_xbar_demux_008:sink_startofpacket
	wire  [58:0] limiter_005_cmd_src_data;                                                                          // limiter_005:cmd_src_data -> cmd_xbar_demux_008:sink_data
	wire   [3:0] limiter_005_cmd_src_channel;                                                                       // limiter_005:cmd_src_channel -> cmd_xbar_demux_008:sink_channel
	wire         limiter_005_cmd_src_ready;                                                                         // cmd_xbar_demux_008:sink_ready -> limiter_005:cmd_src_ready
	wire         rsp_xbar_mux_008_src_endofpacket;                                                                  // rsp_xbar_mux_008:src_endofpacket -> limiter_005:rsp_sink_endofpacket
	wire         rsp_xbar_mux_008_src_valid;                                                                        // rsp_xbar_mux_008:src_valid -> limiter_005:rsp_sink_valid
	wire         rsp_xbar_mux_008_src_startofpacket;                                                                // rsp_xbar_mux_008:src_startofpacket -> limiter_005:rsp_sink_startofpacket
	wire  [58:0] rsp_xbar_mux_008_src_data;                                                                         // rsp_xbar_mux_008:src_data -> limiter_005:rsp_sink_data
	wire   [3:0] rsp_xbar_mux_008_src_channel;                                                                      // rsp_xbar_mux_008:src_channel -> limiter_005:rsp_sink_channel
	wire         rsp_xbar_mux_008_src_ready;                                                                        // limiter_005:rsp_sink_ready -> rsp_xbar_mux_008:src_ready
	wire         cmd_xbar_demux_008_src0_ready;                                                                     // led_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src0_ready
	wire         id_router_013_src_endofpacket;                                                                     // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire         id_router_013_src_valid;                                                                           // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire         id_router_013_src_startofpacket;                                                                   // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [58:0] id_router_013_src_data;                                                                            // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [3:0] id_router_013_src_channel;                                                                         // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire         id_router_013_src_ready;                                                                           // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire         cmd_xbar_demux_008_src1_ready;                                                                     // sw_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src1_ready
	wire         id_router_014_src_endofpacket;                                                                     // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire         id_router_014_src_valid;                                                                           // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire         id_router_014_src_startofpacket;                                                                   // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [58:0] id_router_014_src_data;                                                                            // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [3:0] id_router_014_src_channel;                                                                         // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire         id_router_014_src_ready;                                                                           // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire         cmd_xbar_demux_008_src2_ready;                                                                     // pb_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src2_ready
	wire         id_router_015_src_endofpacket;                                                                     // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire         id_router_015_src_valid;                                                                           // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire         id_router_015_src_startofpacket;                                                                   // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [58:0] id_router_015_src_data;                                                                            // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [3:0] id_router_015_src_channel;                                                                         // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire         id_router_015_src_ready;                                                                           // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire         cmd_xbar_demux_008_src3_ready;                                                                     // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src3_ready
	wire         id_router_016_src_endofpacket;                                                                     // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire         id_router_016_src_valid;                                                                           // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire         id_router_016_src_startofpacket;                                                                   // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [58:0] id_router_016_src_data;                                                                            // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [3:0] id_router_016_src_channel;                                                                         // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire         id_router_016_src_ready;                                                                           // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                  // cmd_xbar_mux_002:src_endofpacket -> width_adapter:in_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                        // cmd_xbar_mux_002:src_valid -> width_adapter:in_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                // cmd_xbar_mux_002:src_startofpacket -> width_adapter:in_startofpacket
	wire  [88:0] cmd_xbar_mux_002_src_data;                                                                         // cmd_xbar_mux_002:src_data -> width_adapter:in_data
	wire  [12:0] cmd_xbar_mux_002_src_channel;                                                                      // cmd_xbar_mux_002:src_channel -> width_adapter:in_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                        // width_adapter:in_ready -> cmd_xbar_mux_002:src_ready
	wire         width_adapter_src_endofpacket;                                                                     // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire         width_adapter_src_valid;                                                                           // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire         width_adapter_src_startofpacket;                                                                   // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [70:0] width_adapter_src_data;                                                                            // width_adapter:out_data -> burst_adapter:sink0_data
	wire         width_adapter_src_ready;                                                                           // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire  [12:0] width_adapter_src_channel;                                                                         // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire         id_router_002_src_endofpacket;                                                                     // id_router_002:src_endofpacket -> width_adapter_001:in_endofpacket
	wire         id_router_002_src_valid;                                                                           // id_router_002:src_valid -> width_adapter_001:in_valid
	wire         id_router_002_src_startofpacket;                                                                   // id_router_002:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [70:0] id_router_002_src_data;                                                                            // id_router_002:src_data -> width_adapter_001:in_data
	wire  [12:0] id_router_002_src_channel;                                                                         // id_router_002:src_channel -> width_adapter_001:in_channel
	wire         id_router_002_src_ready;                                                                           // width_adapter_001:in_ready -> id_router_002:src_ready
	wire         width_adapter_001_src_endofpacket;                                                                 // width_adapter_001:out_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         width_adapter_001_src_valid;                                                                       // width_adapter_001:out_valid -> rsp_xbar_demux_002:sink_valid
	wire         width_adapter_001_src_startofpacket;                                                               // width_adapter_001:out_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [88:0] width_adapter_001_src_data;                                                                        // width_adapter_001:out_data -> rsp_xbar_demux_002:sink_data
	wire         width_adapter_001_src_ready;                                                                       // rsp_xbar_demux_002:sink_ready -> width_adapter_001:out_ready
	wire  [12:0] width_adapter_001_src_channel;                                                                     // width_adapter_001:out_channel -> rsp_xbar_demux_002:sink_channel
	wire         crosser_out_endofpacket;                                                                           // crosser:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         crosser_out_valid;                                                                                 // crosser:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         crosser_out_startofpacket;                                                                         // crosser:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] crosser_out_data;                                                                                  // crosser:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] crosser_out_channel;                                                                               // crosser:out_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                               // cmd_xbar_demux_001:src3_endofpacket -> crosser:in_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                     // cmd_xbar_demux_001:src3_valid -> crosser:in_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                             // cmd_xbar_demux_001:src3_startofpacket -> crosser:in_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src3_data;                                                                      // cmd_xbar_demux_001:src3_data -> crosser:in_data
	wire  [12:0] cmd_xbar_demux_001_src3_channel;                                                                   // cmd_xbar_demux_001:src3_channel -> crosser:in_channel
	wire         cmd_xbar_demux_001_src3_ready;                                                                     // crosser:in_ready -> cmd_xbar_demux_001:src3_ready
	wire         crosser_001_out_endofpacket;                                                                       // crosser_001:out_endofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         crosser_001_out_valid;                                                                             // crosser_001:out_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         crosser_001_out_startofpacket;                                                                     // crosser_001:out_startofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] crosser_001_out_data;                                                                              // crosser_001:out_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] crosser_001_out_channel;                                                                           // crosser_001:out_channel -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                               // cmd_xbar_demux_001:src5_endofpacket -> crosser_001:in_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                     // cmd_xbar_demux_001:src5_valid -> crosser_001:in_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                             // cmd_xbar_demux_001:src5_startofpacket -> crosser_001:in_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src5_data;                                                                      // cmd_xbar_demux_001:src5_data -> crosser_001:in_data
	wire  [12:0] cmd_xbar_demux_001_src5_channel;                                                                   // cmd_xbar_demux_001:src5_channel -> crosser_001:in_channel
	wire         cmd_xbar_demux_001_src5_ready;                                                                     // crosser_001:in_ready -> cmd_xbar_demux_001:src5_ready
	wire         crosser_002_out_endofpacket;                                                                       // crosser_002:out_endofpacket -> sys_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         crosser_002_out_valid;                                                                             // crosser_002:out_valid -> sys_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         crosser_002_out_startofpacket;                                                                     // crosser_002:out_startofpacket -> sys_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] crosser_002_out_data;                                                                              // crosser_002:out_data -> sys_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] crosser_002_out_channel;                                                                           // crosser_002:out_channel -> sys_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                               // cmd_xbar_demux_001:src6_endofpacket -> crosser_002:in_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                     // cmd_xbar_demux_001:src6_valid -> crosser_002:in_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                             // cmd_xbar_demux_001:src6_startofpacket -> crosser_002:in_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src6_data;                                                                      // cmd_xbar_demux_001:src6_data -> crosser_002:in_data
	wire  [12:0] cmd_xbar_demux_001_src6_channel;                                                                   // cmd_xbar_demux_001:src6_channel -> crosser_002:in_channel
	wire         cmd_xbar_demux_001_src6_ready;                                                                     // crosser_002:in_ready -> cmd_xbar_demux_001:src6_ready
	wire         crosser_003_out_endofpacket;                                                                       // crosser_003:out_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         crosser_003_out_valid;                                                                             // crosser_003:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         crosser_003_out_startofpacket;                                                                     // crosser_003:out_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] crosser_003_out_data;                                                                              // crosser_003:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [12:0] crosser_003_out_channel;                                                                           // crosser_003:out_channel -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src12_endofpacket;                                                              // cmd_xbar_demux_001:src12_endofpacket -> crosser_003:in_endofpacket
	wire         cmd_xbar_demux_001_src12_valid;                                                                    // cmd_xbar_demux_001:src12_valid -> crosser_003:in_valid
	wire         cmd_xbar_demux_001_src12_startofpacket;                                                            // cmd_xbar_demux_001:src12_startofpacket -> crosser_003:in_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src12_data;                                                                     // cmd_xbar_demux_001:src12_data -> crosser_003:in_data
	wire  [12:0] cmd_xbar_demux_001_src12_channel;                                                                  // cmd_xbar_demux_001:src12_channel -> crosser_003:in_channel
	wire         cmd_xbar_demux_001_src12_ready;                                                                    // crosser_003:in_ready -> cmd_xbar_demux_001:src12_ready
	wire         crosser_004_out_endofpacket;                                                                       // crosser_004:out_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         crosser_004_out_valid;                                                                             // crosser_004:out_valid -> rsp_xbar_mux_001:sink3_valid
	wire         crosser_004_out_startofpacket;                                                                     // crosser_004:out_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [88:0] crosser_004_out_data;                                                                              // crosser_004:out_data -> rsp_xbar_mux_001:sink3_data
	wire  [12:0] crosser_004_out_channel;                                                                           // crosser_004:out_channel -> rsp_xbar_mux_001:sink3_channel
	wire         crosser_004_out_ready;                                                                             // rsp_xbar_mux_001:sink3_ready -> crosser_004:out_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                               // rsp_xbar_demux_003:src0_endofpacket -> crosser_004:in_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                     // rsp_xbar_demux_003:src0_valid -> crosser_004:in_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                             // rsp_xbar_demux_003:src0_startofpacket -> crosser_004:in_startofpacket
	wire  [88:0] rsp_xbar_demux_003_src0_data;                                                                      // rsp_xbar_demux_003:src0_data -> crosser_004:in_data
	wire  [12:0] rsp_xbar_demux_003_src0_channel;                                                                   // rsp_xbar_demux_003:src0_channel -> crosser_004:in_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                     // crosser_004:in_ready -> rsp_xbar_demux_003:src0_ready
	wire         crosser_005_out_endofpacket;                                                                       // crosser_005:out_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         crosser_005_out_valid;                                                                             // crosser_005:out_valid -> rsp_xbar_mux_001:sink5_valid
	wire         crosser_005_out_startofpacket;                                                                     // crosser_005:out_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [88:0] crosser_005_out_data;                                                                              // crosser_005:out_data -> rsp_xbar_mux_001:sink5_data
	wire  [12:0] crosser_005_out_channel;                                                                           // crosser_005:out_channel -> rsp_xbar_mux_001:sink5_channel
	wire         crosser_005_out_ready;                                                                             // rsp_xbar_mux_001:sink5_ready -> crosser_005:out_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                               // rsp_xbar_demux_005:src0_endofpacket -> crosser_005:in_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                     // rsp_xbar_demux_005:src0_valid -> crosser_005:in_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                             // rsp_xbar_demux_005:src0_startofpacket -> crosser_005:in_startofpacket
	wire  [88:0] rsp_xbar_demux_005_src0_data;                                                                      // rsp_xbar_demux_005:src0_data -> crosser_005:in_data
	wire  [12:0] rsp_xbar_demux_005_src0_channel;                                                                   // rsp_xbar_demux_005:src0_channel -> crosser_005:in_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                     // crosser_005:in_ready -> rsp_xbar_demux_005:src0_ready
	wire         crosser_006_out_endofpacket;                                                                       // crosser_006:out_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         crosser_006_out_valid;                                                                             // crosser_006:out_valid -> rsp_xbar_mux_001:sink6_valid
	wire         crosser_006_out_startofpacket;                                                                     // crosser_006:out_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [88:0] crosser_006_out_data;                                                                              // crosser_006:out_data -> rsp_xbar_mux_001:sink6_data
	wire  [12:0] crosser_006_out_channel;                                                                           // crosser_006:out_channel -> rsp_xbar_mux_001:sink6_channel
	wire         crosser_006_out_ready;                                                                             // rsp_xbar_mux_001:sink6_ready -> crosser_006:out_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                               // rsp_xbar_demux_006:src0_endofpacket -> crosser_006:in_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                     // rsp_xbar_demux_006:src0_valid -> crosser_006:in_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                             // rsp_xbar_demux_006:src0_startofpacket -> crosser_006:in_startofpacket
	wire  [88:0] rsp_xbar_demux_006_src0_data;                                                                      // rsp_xbar_demux_006:src0_data -> crosser_006:in_data
	wire  [12:0] rsp_xbar_demux_006_src0_channel;                                                                   // rsp_xbar_demux_006:src0_channel -> crosser_006:in_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                     // crosser_006:in_ready -> rsp_xbar_demux_006:src0_ready
	wire         crosser_007_out_endofpacket;                                                                       // crosser_007:out_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire         crosser_007_out_valid;                                                                             // crosser_007:out_valid -> rsp_xbar_mux_001:sink12_valid
	wire         crosser_007_out_startofpacket;                                                                     // crosser_007:out_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [88:0] crosser_007_out_data;                                                                              // crosser_007:out_data -> rsp_xbar_mux_001:sink12_data
	wire  [12:0] crosser_007_out_channel;                                                                           // crosser_007:out_channel -> rsp_xbar_mux_001:sink12_channel
	wire         crosser_007_out_ready;                                                                             // rsp_xbar_mux_001:sink12_ready -> crosser_007:out_ready
	wire         rsp_xbar_demux_012_src0_endofpacket;                                                               // rsp_xbar_demux_012:src0_endofpacket -> crosser_007:in_endofpacket
	wire         rsp_xbar_demux_012_src0_valid;                                                                     // rsp_xbar_demux_012:src0_valid -> crosser_007:in_valid
	wire         rsp_xbar_demux_012_src0_startofpacket;                                                             // rsp_xbar_demux_012:src0_startofpacket -> crosser_007:in_startofpacket
	wire  [88:0] rsp_xbar_demux_012_src0_data;                                                                      // rsp_xbar_demux_012:src0_data -> crosser_007:in_data
	wire  [12:0] rsp_xbar_demux_012_src0_channel;                                                                   // rsp_xbar_demux_012:src0_channel -> crosser_007:in_channel
	wire         rsp_xbar_demux_012_src0_ready;                                                                     // crosser_007:in_ready -> rsp_xbar_demux_012:src0_ready
	wire  [12:0] limiter_cmd_valid_data;                                                                            // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire  [12:0] limiter_001_cmd_valid_data;                                                                        // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire  [12:0] limiter_002_cmd_valid_data;                                                                        // limiter_002:cmd_src_valid -> cmd_xbar_demux_002:sink_valid
	wire  [12:0] limiter_003_cmd_valid_data;                                                                        // limiter_003:cmd_src_valid -> cmd_xbar_demux_004:sink_valid
	wire  [12:0] limiter_004_cmd_valid_data;                                                                        // limiter_004:cmd_src_valid -> cmd_xbar_demux_007:sink_valid
	wire   [3:0] limiter_005_cmd_valid_data;                                                                        // limiter_005:cmd_src_valid -> cmd_xbar_demux_008:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                          // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver3_irq;                                                                          // sgdma_tx:csr_irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                                          // sgdma_rx:csr_irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu_d_irq_irq;                                                                                     // irq_mapper:sender_irq -> cpu:d_irq
	wire         irq_mapper_receiver1_irq;                                                                          // irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                                                     // high_res_timer:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver2_irq;                                                                          // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                                                 // sys_timer:irq -> irq_synchronizer_001:receiver_irq

	DE4_SOPC_onchip_memory onchip_memory (
		.clk        (pll_sys_clk),                                                //   clk1.clk
		.address    (onchip_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (onchip_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (onchip_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (onchip_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (onchip_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (onchip_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                              // reset1.reset
	);

	DE4_SOPC_jtag_uart jtag_uart (
		.clk            (pll_sys_clk),                                                            //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.dataavailable  (),                                                                       //                  .dataavailable
		.readyfordata   (),                                                                       //                  .readyfordata
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	DE4_SOPC_high_res_timer high_res_timer (
		.clk        (pll_peripheral_clk),                                          //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                         // reset.reset_n
		.address    (high_res_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (high_res_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (high_res_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (high_res_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~high_res_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)                                //   irq.irq
	);

	DE4_SOPC_sys_timer sys_timer (
		.clk        (pll_peripheral_clk),                                     //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    // reset.reset_n
		.address    (sys_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (sys_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (sys_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (sys_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~sys_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)                       //   irq.irq
	);

	DE4_SOPC_tse_mac tse_mac (
		.ff_tx_data     (sgdma_tx_out_data),                                               //                      transmit.data
		.ff_tx_eop      (sgdma_tx_out_endofpacket),                                        //                              .endofpacket
		.ff_tx_err      (sgdma_tx_out_error),                                              //                              .error
		.ff_tx_mod      (sgdma_tx_out_empty),                                              //                              .empty
		.ff_tx_rdy      (sgdma_tx_out_ready),                                              //                              .ready
		.ff_tx_sop      (sgdma_tx_out_startofpacket),                                      //                              .startofpacket
		.ff_tx_wren     (sgdma_tx_out_valid),                                              //                              .valid
		.ff_tx_clk      (pll_sys_clk),                                                     //      receive_clock_connection.clk
		.ff_rx_data     (tse_mac_receive_data),                                            //                       receive.data
		.ff_rx_dval     (tse_mac_receive_valid),                                           //                              .valid
		.ff_rx_eop      (tse_mac_receive_endofpacket),                                     //                              .endofpacket
		.ff_rx_mod      (tse_mac_receive_empty),                                           //                              .empty
		.ff_rx_rdy      (tse_mac_receive_ready),                                           //                              .ready
		.ff_rx_sop      (tse_mac_receive_startofpacket),                                   //                              .startofpacket
		.rx_err         (tse_mac_receive_error),                                           //                              .error
		.ff_rx_clk      (pll_sys_clk),                                                     //     transmit_clock_connection.clk
		.address        (tse_mac_control_port_translator_avalon_anti_slave_0_address),     //                  control_port.address
		.readdata       (tse_mac_control_port_translator_avalon_anti_slave_0_readdata),    //                              .readdata
		.read           (tse_mac_control_port_translator_avalon_anti_slave_0_read),        //                              .read
		.writedata      (tse_mac_control_port_translator_avalon_anti_slave_0_writedata),   //                              .writedata
		.write          (tse_mac_control_port_translator_avalon_anti_slave_0_write),       //                              .write
		.waitrequest    (tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest), //                              .waitrequest
		.clk            (pll_sys_clk),                                                     // control_port_clock_connection.clk
		.reset          (rst_controller_reset_out_reset),                                  //              reset_connection.reset
		.mdio_out       (mdio_out_from_the_tse_mac),                                       //            conduit_connection.export
		.mdio_oen       (mdio_oen_from_the_tse_mac),                                       //                              .export
		.mdio_in        (mdio_in_to_the_tse_mac),                                          //                              .export
		.mdc            (mdc_from_the_tse_mac),                                            //                              .export
		.led_an         (led_an_from_the_tse_mac),                                         //                              .export
		.led_char_err   (led_char_err_from_the_tse_mac),                                   //                              .export
		.led_link       (led_link_from_the_tse_mac),                                       //                              .export
		.led_disp_err   (led_disp_err_from_the_tse_mac),                                   //                              .export
		.led_crs        (led_crs_from_the_tse_mac),                                        //                              .export
		.led_col        (led_col_from_the_tse_mac),                                        //                              .export
		.txp            (txp_from_the_tse_mac),                                            //                              .export
		.rxp            (rxp_to_the_tse_mac),                                              //                              .export
		.ref_clk        (ref_clk_to_the_tse_mac),                                          //                              .export
		.rx_recovclkout (rx_recovclkout_from_the_tse_mac)                                  //                              .export
	);

	DE4_SOPC_sgdma_tx sgdma_tx (
		.clk                           (pll_sys_clk),                                            //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),                        //            reset.reset_n
		.csr_chipselect                (sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect), //              csr.chipselect
		.csr_address                   (sgdma_tx_csr_translator_avalon_anti_slave_0_address),    //                 .address
		.csr_read                      (sgdma_tx_csr_translator_avalon_anti_slave_0_read),       //                 .read
		.csr_write                     (sgdma_tx_csr_translator_avalon_anti_slave_0_write),      //                 .write
		.csr_writedata                 (sgdma_tx_csr_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.csr_readdata                  (sgdma_tx_csr_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),                      //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),                 //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),                   //                 .waitrequest
		.descriptor_read_address       (sgdma_tx_descriptor_read_address),                       //                 .address
		.descriptor_read_read          (sgdma_tx_descriptor_read_read),                          //                 .read
		.descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),                  // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_tx_descriptor_write_address),                      //                 .address
		.descriptor_write_write        (sgdma_tx_descriptor_write_write),                        //                 .write
		.descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),                    //                 .writedata
		.csr_irq                       (irq_mapper_receiver3_irq),                               //          csr_irq.irq
		.m_read_readdata               (sgdma_tx_m_read_readdata),                               //           m_read.readdata
		.m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),                          //                 .readdatavalid
		.m_read_waitrequest            (sgdma_tx_m_read_waitrequest),                            //                 .waitrequest
		.m_read_address                (sgdma_tx_m_read_address),                                //                 .address
		.m_read_read                   (sgdma_tx_m_read_read),                                   //                 .read
		.out_data                      (sgdma_tx_out_data),                                      //              out.data
		.out_valid                     (sgdma_tx_out_valid),                                     //                 .valid
		.out_ready                     (sgdma_tx_out_ready),                                     //                 .ready
		.out_endofpacket               (sgdma_tx_out_endofpacket),                               //                 .endofpacket
		.out_startofpacket             (sgdma_tx_out_startofpacket),                             //                 .startofpacket
		.out_empty                     (sgdma_tx_out_empty),                                     //                 .empty
		.out_error                     (sgdma_tx_out_error)                                      //                 .error
	);

	DE4_SOPC_sgdma_rx sgdma_rx (
		.clk                           (pll_sys_clk),                                            //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),                        //            reset.reset_n
		.csr_chipselect                (sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect), //              csr.chipselect
		.csr_address                   (sgdma_rx_csr_translator_avalon_anti_slave_0_address),    //                 .address
		.csr_read                      (sgdma_rx_csr_translator_avalon_anti_slave_0_read),       //                 .read
		.csr_write                     (sgdma_rx_csr_translator_avalon_anti_slave_0_write),      //                 .write
		.csr_writedata                 (sgdma_rx_csr_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.csr_readdata                  (sgdma_rx_csr_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),                      //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),                 //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),                   //                 .waitrequest
		.descriptor_read_address       (sgdma_rx_descriptor_read_address),                       //                 .address
		.descriptor_read_read          (sgdma_rx_descriptor_read_read),                          //                 .read
		.descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),                  // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_rx_descriptor_write_address),                      //                 .address
		.descriptor_write_write        (sgdma_rx_descriptor_write_write),                        //                 .write
		.descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),                    //                 .writedata
		.csr_irq                       (irq_mapper_receiver4_irq),                               //          csr_irq.irq
		.m_write_waitrequest           (sgdma_rx_m_write_waitrequest),                           //          m_write.waitrequest
		.m_write_address               (sgdma_rx_m_write_address),                               //                 .address
		.m_write_write                 (sgdma_rx_m_write_write),                                 //                 .write
		.m_write_writedata             (sgdma_rx_m_write_writedata),                             //                 .writedata
		.m_write_byteenable            (sgdma_rx_m_write_byteenable),                            //                 .byteenable
		.in_startofpacket              (tse_mac_receive_startofpacket),                          //               in.startofpacket
		.in_endofpacket                (tse_mac_receive_endofpacket),                            //                 .endofpacket
		.in_empty                      (tse_mac_receive_empty),                                  //                 .empty
		.in_data                       (tse_mac_receive_data),                                   //                 .data
		.in_valid                      (tse_mac_receive_valid),                                  //                 .valid
		.in_ready                      (tse_mac_receive_ready),                                  //                 .ready
		.in_error                      (tse_mac_receive_error)                                   //                 .error
	);

	DE4_SOPC_descriptor_memory descriptor_memory (
		.clk        (pll_sys_clk),                                                    //   clk1.clk
		.address    (descriptor_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (descriptor_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (descriptor_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (descriptor_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (descriptor_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                                  // reset1.reset
	);

	DE4_SOPC_led_pio led_pio (
		.clk        (pll_peripheral_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address    (led_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_port_from_the_led_pio)                             // external_connection.export
	);

	DE4_SOPC_sw_pio sw_pio (
		.clk      (pll_peripheral_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),               //               reset.reset_n
		.address  (sw_pio_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (sw_pio_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (in_port_to_the_sw_pio)                              // external_connection.export
	);

	DE4_SOPC_pb_pio pb_pio (
		.clk      (pll_peripheral_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),               //               reset.reset_n
		.address  (pb_pio_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (pb_pio_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (in_port_to_the_pb_pio)                              // external_connection.export
	);

	DE4_SOPC_seven_seg_pio seven_seg_pio (
		.clk        (pll_peripheral_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                        //               reset.reset_n
		.address    (seven_seg_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~seven_seg_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (seven_seg_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (seven_seg_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (seven_seg_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_port_from_the_seven_seg_pio)                             // external_connection.export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (6),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) peripheral_clock_crossing (
		.m0_clk           (pll_peripheral_clk),                                                        //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                                        // m0_reset.reset
		.s0_clk           (pll_sys_clk),                                                               //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                                            // s0_reset.reset
		.s0_waitrequest   (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (peripheral_clock_crossing_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (peripheral_clock_crossing_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (peripheral_clock_crossing_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (peripheral_clock_crossing_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (peripheral_clock_crossing_m0_writedata),                                    //         .writedata
		.m0_address       (peripheral_clock_crossing_m0_address),                                      //         .address
		.m0_write         (peripheral_clock_crossing_m0_write),                                        //         .write
		.m0_read          (peripheral_clock_crossing_m0_read),                                         //         .read
		.m0_byteenable    (peripheral_clock_crossing_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (peripheral_clock_crossing_m0_debugaccess)                                   //         .debugaccess
	);

	DE4_SOPC_cpu cpu (
		.clk                                   (pll_sys_clk),                                                        //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                    //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                          //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                                      //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	DE4_SOPC_sysid sysid (
		.clock    (pll_peripheral_clk),                                          //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                         //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	DE4_SOPC_flash_tristate_bridge_bridge_0 flash_tristate_bridge_bridge_0 (
		.clk                                  (pll_sys_clk),                                                             //   clk.clk
		.reset                                (rst_controller_reset_out_reset),                                          // reset.reset
		.request                              (flash_tristate_bridge_pinsharer_0_tcm_request),                           //   tcs.request
		.grant                                (flash_tristate_bridge_pinsharer_0_tcm_grant),                             //      .grant
		.tcs_flash_tristate_bridge_address    (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_address_out), //      .flash_tristate_bridge_address_out
		.tcs_flash_tristate_bridge_writen     (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_writen_out),  //      .flash_tristate_bridge_writen_out
		.tcs_flash_tristate_bridge_data       (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_out),    //      .flash_tristate_bridge_data_out
		.tcs_flash_tristate_bridge_data_outen (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_outen),  //      .flash_tristate_bridge_data_outen
		.tcs_flash_tristate_bridge_data_in    (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_in),     //      .flash_tristate_bridge_data_in
		.tcs_select_n_to_the_ext_flash        (flash_tristate_bridge_pinsharer_0_tcm_select_n_to_the_ext_flash_out),     //      .select_n_to_the_ext_flash_out
		.tcs_flash_tristate_bridge_readn      (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_readn_out),   //      .flash_tristate_bridge_readn_out
		.flash_tristate_bridge_address        (flash_tristate_bridge_address),                                           //   out.flash_tristate_bridge_address
		.flash_tristate_bridge_writen         (flash_tristate_bridge_writen),                                            //      .flash_tristate_bridge_writen
		.flash_tristate_bridge_data           (flash_tristate_bridge_data),                                              //      .flash_tristate_bridge_data
		.select_n_to_the_ext_flash            (select_n_to_the_ext_flash),                                               //      .select_n_to_the_ext_flash
		.flash_tristate_bridge_readn          (flash_tristate_bridge_readn)                                              //      .flash_tristate_bridge_readn
	);

	DE4_SOPC_flash_tristate_bridge_pinSharer_0 flash_tristate_bridge_pinsharer_0 (
		.clk_clk                          (pll_sys_clk),                                                             //   clk.clk
		.reset_reset                      (rst_controller_reset_out_reset),                                          // reset.reset
		.request                          (flash_tristate_bridge_pinsharer_0_tcm_request),                           //   tcm.request
		.grant                            (flash_tristate_bridge_pinsharer_0_tcm_grant),                             //      .grant
		.flash_tristate_bridge_address    (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_address_out), //      .flash_tristate_bridge_address_out
		.flash_tristate_bridge_readn      (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_readn_out),   //      .flash_tristate_bridge_readn_out
		.flash_tristate_bridge_writen     (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_writen_out),  //      .flash_tristate_bridge_writen_out
		.flash_tristate_bridge_data       (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_out),    //      .flash_tristate_bridge_data_out
		.flash_tristate_bridge_data_in    (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_in),     //      .flash_tristate_bridge_data_in
		.flash_tristate_bridge_data_outen (flash_tristate_bridge_pinsharer_0_tcm_flash_tristate_bridge_data_outen),  //      .flash_tristate_bridge_data_outen
		.select_n_to_the_ext_flash        (flash_tristate_bridge_pinsharer_0_tcm_select_n_to_the_ext_flash_out),     //      .select_n_to_the_ext_flash_out
		.tcs0_request                     (ext_flash_tcm_request),                                                   //  tcs0.request
		.tcs0_grant                       (ext_flash_tcm_grant),                                                     //      .grant
		.tcs0_address_out                 (ext_flash_tcm_address_out),                                               //      .address_out
		.tcs0_read_n_out                  (ext_flash_tcm_read_n_out),                                                //      .read_n_out
		.tcs0_write_n_out                 (ext_flash_tcm_write_n_out),                                               //      .write_n_out
		.tcs0_data_out                    (ext_flash_tcm_data_out),                                                  //      .data_out
		.tcs0_data_in                     (ext_flash_tcm_data_in),                                                   //      .data_in
		.tcs0_data_outen                  (ext_flash_tcm_data_outen),                                                //      .data_outen
		.tcs0_chipselect_n_out            (ext_flash_tcm_chipselect_n_out)                                           //      .chipselect_n_out
	);

	DE4_SOPC_ext_flash #(
		.TCM_ADDRESS_W                  (25),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (100),
		.TCM_WRITE_WAIT                 (100),
		.TCM_SETUP_WAIT                 (25),
		.TCM_DATA_HOLD                  (20),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) ext_flash (
		.clk_clk              (pll_sys_clk),                                                //   clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                             // reset.reset
		.uas_address          (ext_flash_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount       (ext_flash_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read             (ext_flash_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write            (ext_flash_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest      (ext_flash_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (ext_flash_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable       (ext_flash_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata         (ext_flash_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata        (ext_flash_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock             (ext_flash_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess      (ext_flash_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (ext_flash_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_read_n_out       (ext_flash_tcm_read_n_out),                                   //      .read_n_out
		.tcm_chipselect_n_out (ext_flash_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_request          (ext_flash_tcm_request),                                      //      .request
		.tcm_grant            (ext_flash_tcm_grant),                                        //      .grant
		.tcm_address_out      (ext_flash_tcm_address_out),                                  //      .address_out
		.tcm_data_out         (ext_flash_tcm_data_out),                                     //      .data_out
		.tcm_data_outen       (ext_flash_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in          (ext_flash_tcm_data_in)                                       //      .data_in
	);

	DE4_SOPC_altpll_0 altpll_0 (
		.clk       (ext_clk),                                                     //       inclk_interface.clk
		.reset     (rst_controller_002_reset_out_reset),                          // inclk_interface_reset.reset
		.read      (altpll_0_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (altpll_0_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (altpll_0_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (pll_sys_clk),                                                 //                    c0.clk
		.c1        (pll_peripheral_clk),                                          //                    c1.clk
		.areset    (altpll_0_areset_conduit_export),                              //        areset_conduit.export
		.locked    (altpll_0_locked_conduit_export),                              //        locked_conduit.export
		.phasedone (altpll_0_phasedone_conduit_export)                            //     phasedone_conduit.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (27),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                   (pll_sys_clk),                                                               //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address           (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                      //               (terminated)
		.av_byteenable         (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                      //               (terminated)
		.av_begintransfer      (1'b0),                                                                      //               (terminated)
		.av_chipselect         (1'b0),                                                                      //               (terminated)
		.av_write              (1'b0),                                                                      //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock               (1'b0),                                                                      //               (terminated)
		.av_debugaccess        (1'b0),                                                                      //               (terminated)
		.uav_clken             (),                                                                          //               (terminated)
		.av_clken              (1'b1)                                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (27),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_data_master_translator (
		.clk                   (pll_sys_clk),                                                        //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address           (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_data_master_read),                                               //                          .read
		.av_readdata           (cpu_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (cpu_data_master_write),                                              //                          .write
		.av_writedata          (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_rx_descriptor_read_translator (
		.clk                   (pll_sys_clk),                                                                 //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_rx_descriptor_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_rx_descriptor_read_waitrequest),                                        //                          .waitrequest
		.av_read               (sgdma_rx_descriptor_read_read),                                               //                          .read
		.av_readdata           (sgdma_rx_descriptor_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (sgdma_rx_descriptor_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_rx_descriptor_write_translator (
		.clk                   (pll_sys_clk),                                                                  //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                     reset.reset
		.uav_address           (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_rx_descriptor_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_rx_descriptor_write_waitrequest),                                        //                          .waitrequest
		.av_write              (sgdma_rx_descriptor_write_write),                                              //                          .write
		.av_writedata          (sgdma_rx_descriptor_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                         //               (terminated)
		.av_byteenable         (4'b1111),                                                                      //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_read               (1'b0),                                                                         //               (terminated)
		.av_readdata           (),                                                                             //               (terminated)
		.av_readdatavalid      (),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.av_debugaccess        (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_tx_descriptor_read_translator (
		.clk                   (pll_sys_clk),                                                                 //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_tx_descriptor_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_tx_descriptor_read_waitrequest),                                        //                          .waitrequest
		.av_read               (sgdma_tx_descriptor_read_read),                                               //                          .read
		.av_readdata           (sgdma_tx_descriptor_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (sgdma_tx_descriptor_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_tx_descriptor_write_translator (
		.clk                   (pll_sys_clk),                                                                  //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                     reset.reset
		.uav_address           (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_tx_descriptor_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_tx_descriptor_write_waitrequest),                                        //                          .waitrequest
		.av_write              (sgdma_tx_descriptor_write_write),                                              //                          .write
		.av_writedata          (sgdma_tx_descriptor_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                         //               (terminated)
		.av_byteenable         (4'b1111),                                                                      //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                         //               (terminated)
		.av_begintransfer      (1'b0),                                                                         //               (terminated)
		.av_chipselect         (1'b0),                                                                         //               (terminated)
		.av_read               (1'b0),                                                                         //               (terminated)
		.av_readdata           (),                                                                             //               (terminated)
		.av_readdatavalid      (),                                                                             //               (terminated)
		.av_lock               (1'b0),                                                                         //               (terminated)
		.av_debugaccess        (1'b0),                                                                         //               (terminated)
		.uav_clken             (),                                                                             //               (terminated)
		.av_clken              (1'b1)                                                                          //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_rx_m_write_translator (
		.clk                   (pll_sys_clk),                                                         //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                      //                     reset.reset
		.uav_address           (sgdma_rx_m_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_rx_m_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_rx_m_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_rx_m_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_rx_m_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_rx_m_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_rx_m_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_rx_m_write_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (sgdma_rx_m_write_byteenable),                                         //                          .byteenable
		.av_write              (sgdma_rx_m_write_write),                                              //                          .write
		.av_writedata          (sgdma_rx_m_write_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                //               (terminated)
		.av_begintransfer      (1'b0),                                                                //               (terminated)
		.av_chipselect         (1'b0),                                                                //               (terminated)
		.av_read               (1'b0),                                                                //               (terminated)
		.av_readdata           (),                                                                    //               (terminated)
		.av_readdatavalid      (),                                                                    //               (terminated)
		.av_lock               (1'b0),                                                                //               (terminated)
		.av_debugaccess        (1'b0),                                                                //               (terminated)
		.uav_clken             (),                                                                    //               (terminated)
		.av_clken              (1'b1)                                                                 //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_tx_m_read_translator (
		.clk                   (pll_sys_clk),                                                        //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address           (sgdma_tx_m_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sgdma_tx_m_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sgdma_tx_m_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sgdma_tx_m_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sgdma_tx_m_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sgdma_tx_m_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sgdma_tx_m_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sgdma_tx_m_read_waitrequest),                                        //                          .waitrequest
		.av_read               (sgdma_tx_m_read_read),                                               //                          .read
		.av_readdata           (sgdma_tx_m_read_readdata),                                           //                          .readdata
		.av_readdatavalid      (sgdma_tx_m_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_byteenable         (4'b1111),                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_write              (1'b0),                                                               //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                               //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                   (pll_sys_clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (17),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory_s1_translator (
		.clk                   (pll_sys_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (onchip_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (onchip_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (onchip_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (onchip_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (onchip_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (onchip_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (onchip_memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (25),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (2),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ext_flash_uas_translator (
		.clk                   (pll_sys_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ext_flash_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ext_flash_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ext_flash_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ext_flash_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ext_flash_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (ext_flash_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (ext_flash_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (ext_flash_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (ext_flash_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock               (ext_flash_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess        (ext_flash_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                   (pll_peripheral_clk),                                                             //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                             //                    reset.reset
		.uav_address           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                               //              (terminated)
		.av_read               (),                                                                               //              (terminated)
		.av_writedata          (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                   (pll_sys_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_byteenable         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) high_res_timer_s1_translator (
		.clk                   (pll_peripheral_clk),                                                           //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (high_res_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (high_res_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (high_res_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (high_res_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (high_res_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sys_timer_s1_translator (
		.clk                   (pll_peripheral_clk),                                                      //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address           (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sys_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sys_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sys_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sys_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sys_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                        //              (terminated)
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) tse_mac_control_port_translator (
		.clk                   (pll_sys_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (tse_mac_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (tse_mac_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (tse_mac_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (tse_mac_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (tse_mac_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_byteenable         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.av_chipselect         (),                                                                                //              (terminated)
		.av_clken              (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sgdma_tx_csr_translator (
		.clk                   (pll_sys_clk),                                                             //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sgdma_tx_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sgdma_tx_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sgdma_tx_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sgdma_tx_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sgdma_tx_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sgdma_rx_csr_translator (
		.clk                   (pll_sys_clk),                                                             //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sgdma_rx_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sgdma_rx_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sgdma_rx_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sgdma_rx_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sgdma_rx_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                        //              (terminated)
		.av_burstcount         (),                                                                        //              (terminated)
		.av_byteenable         (),                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                        //              (terminated)
		.av_lock               (),                                                                        //              (terminated)
		.av_clken              (),                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                    //              (terminated)
		.av_debugaccess        (),                                                                        //              (terminated)
		.av_outputenable       ()                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) descriptor_memory_s1_translator (
		.clk                   (pll_sys_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (descriptor_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (descriptor_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (descriptor_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (descriptor_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (descriptor_memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                                //              (terminated)
		.av_begintransfer      (),                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                //              (terminated)
		.av_burstcount         (),                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                //              (terminated)
		.av_lock               (),                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                //              (terminated)
		.av_outputenable       ()                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (6),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) peripheral_clock_crossing_s0_translator (
		.clk                   (pll_sys_clk),                                                                             //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                          //                    reset.reset
		.uav_address           (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (peripheral_clock_crossing_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                                        //              (terminated)
		.av_lock               (),                                                                                        //              (terminated)
		.av_chipselect         (),                                                                                        //              (terminated)
		.av_clken              (),                                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) altpll_0_pll_slave_translator (
		.clk                   (ext_clk),                                                                       //                      clk.clk
		.reset                 (rst_controller_002_reset_out_reset),                                            //                    reset.reset
		.uav_address           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (altpll_0_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (altpll_0_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (altpll_0_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_waitrequest        (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (6),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (6),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) peripheral_clock_crossing_m0_translator (
		.clk                   (pll_peripheral_clk),                                                              //                       clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                              //                     reset.reset
		.uav_address           (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (peripheral_clock_crossing_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (peripheral_clock_crossing_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (peripheral_clock_crossing_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (peripheral_clock_crossing_m0_byteenable),                                         //                          .byteenable
		.av_read               (peripheral_clock_crossing_m0_read),                                               //                          .read
		.av_readdata           (peripheral_clock_crossing_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (peripheral_clock_crossing_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (peripheral_clock_crossing_m0_write),                                              //                          .write
		.av_writedata          (peripheral_clock_crossing_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (peripheral_clock_crossing_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                                            //               (terminated)
		.av_begintransfer      (1'b0),                                                                            //               (terminated)
		.av_chipselect         (1'b0),                                                                            //               (terminated)
		.av_lock               (1'b0),                                                                            //               (terminated)
		.uav_clken             (),                                                                                //               (terminated)
		.av_clken              (1'b1)                                                                             //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (6),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_pio_s1_translator (
		.clk                   (pll_peripheral_clk),                                                    //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (led_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (led_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (led_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (led_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (led_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (6),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sw_pio_s1_translator (
		.clk                   (pll_peripheral_clk),                                                   //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address           (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sw_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sw_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_writedata          (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (6),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pb_pio_s1_translator (
		.clk                   (pll_peripheral_clk),                                                   //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address           (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pb_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (pb_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_writedata          (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (6),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) seven_seg_pio_s1_translator (
		.clk                   (pll_peripheral_clk),                                                          //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address           (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (seven_seg_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (seven_seg_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (seven_seg_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (seven_seg_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (seven_seg_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) high_res_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_peripheral_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_001_out_ready),                                                                  //              cp.ready
		.cp_valid                (crosser_001_out_valid),                                                                  //                .valid
		.cp_data                 (crosser_001_out_data),                                                                   //                .data
		.cp_startofpacket        (crosser_001_out_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (crosser_001_out_endofpacket),                                                            //                .endofpacket
		.cp_channel              (crosser_001_out_channel),                                                                //                .channel
		.rf_sink_ready           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_peripheral_clk),                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_peripheral_clk),                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_startofpacket  (1'b0),                                                                             // (terminated)
		.in_endofpacket    (1'b0),                                                                             // (terminated)
		.out_startofpacket (),                                                                                 // (terminated)
		.out_endofpacket   (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                   //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (61),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (65),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (69),
		.PKT_DEST_ID_L             (66),
		.PKT_BURSTWRAP_H           (60),
		.PKT_BURSTWRAP_L           (58),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (55),
		.PKT_PROTECTION_H          (70),
		.PKT_PROTECTION_L          (70),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (71),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ext_flash_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                      //                .channel
		.rf_sink_ready           (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (72),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_clk),                                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                    //       clk_reset.reset
		.m0_address              (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                                  //                .channel
		.rf_sink_ready           (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (81),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_clk),                                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.in_data           (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (13),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (6),
		.BURSTWRAP_VALUE           (7)
	) sgdma_rx_m_write_translator_avalon_universal_master_0_agent (
		.clk              (pll_sys_clk),                                                                  //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.av_address       (sgdma_rx_m_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_rx_m_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_rx_m_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_rx_m_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_rx_m_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_rx_m_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_001_src2_valid),                                                //        rp.valid
		.rp_data          (rsp_xbar_demux_001_src2_data),                                                 //          .data
		.rp_channel       (rsp_xbar_demux_001_src2_channel),                                              //          .channel
		.rp_startofpacket (rsp_xbar_demux_001_src2_startofpacket),                                        //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),                                          //          .endofpacket
		.rp_ready         (rsp_xbar_demux_001_src2_ready)                                                 //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sys_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_peripheral_clk),                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sys_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_002_out_ready),                                                             //              cp.ready
		.cp_valid                (crosser_002_out_valid),                                                             //                .valid
		.cp_data                 (crosser_002_out_data),                                                              //                .data
		.cp_startofpacket        (crosser_002_out_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (crosser_002_out_endofpacket),                                                       //                .endofpacket
		.cp_channel              (crosser_002_out_channel),                                                           //                .channel
		.rf_sink_ready           (sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_peripheral_clk),                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sys_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sys_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_peripheral_clk),                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sys_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_startofpacket  (1'b0),                                                                        // (terminated)
		.in_endofpacket    (1'b0),                                                                        // (terminated)
		.out_startofpacket (),                                                                            // (terminated)
		.out_endofpacket   (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (13),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (7)
	) sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent (
		.clk              (pll_sys_clk),                                                                           //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.av_address       (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_010_src2_valid),                                                         //        rp.valid
		.rp_data          (rsp_xbar_demux_010_src2_data),                                                          //          .data
		.rp_channel       (rsp_xbar_demux_010_src2_channel),                                                       //          .channel
		.rp_startofpacket (rsp_xbar_demux_010_src2_startofpacket),                                                 //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_010_src2_endofpacket),                                                   //          .endofpacket
		.rp_ready         (rsp_xbar_demux_010_src2_ready)                                                          //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (13),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (7),
		.BURSTWRAP_VALUE           (7)
	) sgdma_tx_m_read_translator_avalon_universal_master_0_agent (
		.clk              (pll_sys_clk),                                                                 //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.av_address       (sgdma_tx_m_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_tx_m_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_tx_m_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_tx_m_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_tx_m_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_tx_m_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_004_rsp_src_valid),                                                   //        rp.valid
		.rp_data          (limiter_004_rsp_src_data),                                                    //          .data
		.rp_channel       (limiter_004_rsp_src_channel),                                                 //          .channel
		.rp_startofpacket (limiter_004_rsp_src_startofpacket),                                           //          .startofpacket
		.rp_endofpacket   (limiter_004_rsp_src_endofpacket),                                             //          .endofpacket
		.rp_ready         (limiter_004_rsp_src_ready)                                                    //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sgdma_tx_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                   //                .channel
		.rf_sink_ready           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_peripheral_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                        //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                        //                .valid
		.cp_data                 (crosser_out_data),                                                                         //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                                //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                                  //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                      //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_peripheral_clk),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_peripheral_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_startofpacket  (1'b0),                                                                               // (terminated)
		.in_endofpacket    (1'b0),                                                                               // (terminated)
		.out_startofpacket (),                                                                                   // (terminated)
		.out_endofpacket   (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (13),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (4),
		.BURSTWRAP_VALUE           (7)
	) sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent (
		.clk              (pll_sys_clk),                                                                          //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_003_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_003_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_003_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_003_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_003_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_003_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (13),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (5),
		.BURSTWRAP_VALUE           (7)
	) sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent (
		.clk              (pll_sys_clk),                                                                           //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.av_address       (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_010_src4_valid),                                                         //        rp.valid
		.rp_data          (rsp_xbar_demux_010_src4_data),                                                          //          .data
		.rp_channel       (rsp_xbar_demux_010_src4_channel),                                                       //          .channel
		.rp_startofpacket (rsp_xbar_demux_010_src4_startofpacket),                                                 //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_010_src4_endofpacket),                                                   //          .endofpacket
		.rp_ready         (rsp_xbar_demux_010_src4_ready)                                                          //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) tse_mac_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                           //                .channel
		.rf_sink_ready           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sgdma_rx_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                                   //                .channel
		.rf_sink_ready           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (13),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (pll_sys_clk),                                                                        //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address       (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                              //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                               //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                            //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                        //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                               //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) onchip_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                          //                .channel
		.rf_sink_ready           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) descriptor_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_010_src_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_mux_010_src_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_mux_010_src_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_mux_010_src_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_010_src_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_mux_010_src_channel),                                                              //                .channel
		.rf_sink_ready           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (ext_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_003_out_ready),                                                                   //              cp.ready
		.cp_valid                (crosser_003_out_valid),                                                                   //                .valid
		.cp_data                 (crosser_003_out_data),                                                                    //                .data
		.cp_startofpacket        (crosser_003_out_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (crosser_003_out_endofpacket),                                                             //                .endofpacket
		.cp_channel              (crosser_003_out_channel),                                                                 //                .channel
		.rf_sink_ready           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (ext_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (ext_clk),                                                                           //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                // clk_reset.reset
		.in_data           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_startofpacket  (1'b0),                                                                              // (terminated)
		.in_endofpacket    (1'b0),                                                                              // (terminated)
		.out_startofpacket (),                                                                                  // (terminated)
		.out_endofpacket   (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (13),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7)
	) sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent (
		.clk              (pll_sys_clk),                                                                          //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_002_rsp_src_valid),                                                            //        rp.valid
		.rp_data          (limiter_002_rsp_src_data),                                                             //          .data
		.rp_channel       (limiter_002_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket (limiter_002_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (limiter_002_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (limiter_002_rsp_src_ready)                                                             //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.ST_CHANNEL_W              (13),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sys_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sys_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (88),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (13),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk              (pll_sys_clk),                                                                 //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.av_address       (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                   //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                    //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                 //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                           //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                             //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                    //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (58),
		.PKT_PROTECTION_L          (58),
		.PKT_BEGIN_BURST           (53),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_ADDR_H                (41),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (42),
		.PKT_TRANS_POSTED          (43),
		.PKT_TRANS_WRITE           (44),
		.PKT_TRANS_READ            (45),
		.PKT_TRANS_LOCK            (46),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (55),
		.PKT_SRC_ID_L              (54),
		.PKT_DEST_ID_H             (57),
		.PKT_DEST_ID_L             (56),
		.ST_DATA_W                 (59),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7)
	) peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent (
		.clk              (pll_peripheral_clk),                                                                       //       clk.clk
		.reset            (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_005_rsp_src_valid),                                                                //        rp.valid
		.rp_data          (limiter_005_rsp_src_data),                                                                 //          .data
		.rp_channel       (limiter_005_rsp_src_channel),                                                              //          .channel
		.rp_startofpacket (limiter_005_rsp_src_startofpacket),                                                        //          .startofpacket
		.rp_endofpacket   (limiter_005_rsp_src_endofpacket),                                                          //          .endofpacket
		.rp_ready         (limiter_005_rsp_src_ready)                                                                 //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (53),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (41),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (42),
		.PKT_TRANS_POSTED          (43),
		.PKT_TRANS_WRITE           (44),
		.PKT_TRANS_READ            (45),
		.PKT_TRANS_LOCK            (46),
		.PKT_SRC_ID_H              (55),
		.PKT_SRC_ID_L              (54),
		.PKT_DEST_ID_H             (57),
		.PKT_DEST_ID_L             (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (58),
		.PKT_PROTECTION_L          (58),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (59),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) seven_seg_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_peripheral_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src3_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src3_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_008_src3_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src3_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src3_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src3_channel),                                                       //                .channel
		.rf_sink_ready           (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (60),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_peripheral_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (53),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (41),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (42),
		.PKT_TRANS_POSTED          (43),
		.PKT_TRANS_WRITE           (44),
		.PKT_TRANS_READ            (45),
		.PKT_TRANS_LOCK            (46),
		.PKT_SRC_ID_H              (55),
		.PKT_SRC_ID_L              (54),
		.PKT_DEST_ID_H             (57),
		.PKT_DEST_ID_L             (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (58),
		.PKT_PROTECTION_L          (58),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (59),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sw_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_peripheral_clk),                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sw_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src1_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src1_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_008_src1_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src1_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src1_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src1_channel),                                                //                .channel
		.rf_sink_ready           (sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (60),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_peripheral_clk),                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (53),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (41),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (42),
		.PKT_TRANS_POSTED          (43),
		.PKT_TRANS_WRITE           (44),
		.PKT_TRANS_READ            (45),
		.PKT_TRANS_LOCK            (46),
		.PKT_SRC_ID_H              (55),
		.PKT_SRC_ID_L              (54),
		.PKT_DEST_ID_H             (57),
		.PKT_DEST_ID_L             (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (58),
		.PKT_PROTECTION_L          (58),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (59),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) led_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_peripheral_clk),                                                              //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src0_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src0_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_008_src0_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src0_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src0_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src0_channel),                                                 //                .channel
		.rf_sink_ready           (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (60),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_peripheral_clk),                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (53),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (41),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (42),
		.PKT_TRANS_POSTED          (43),
		.PKT_TRANS_WRITE           (44),
		.PKT_TRANS_READ            (45),
		.PKT_TRANS_LOCK            (46),
		.PKT_SRC_ID_H              (55),
		.PKT_SRC_ID_L              (54),
		.PKT_DEST_ID_H             (57),
		.PKT_DEST_ID_L             (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (58),
		.PKT_PROTECTION_L          (58),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (59),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pb_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_peripheral_clk),                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pb_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src2_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src2_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_008_src2_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src2_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src2_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src2_channel),                                                //                .channel
		.rf_sink_ready           (pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pb_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pb_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pb_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pb_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pb_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pb_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (60),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_peripheral_clk),                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pb_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pb_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	DE4_SOPC_addr_router addr_router (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                              //          .valid
		.src_data           (addr_router_src_data),                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                         //          .endofpacket
	);

	DE4_SOPC_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                   //          .valid
		.src_data           (addr_router_001_src_data),                                                    //          .data
		.src_channel        (addr_router_001_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                              //          .endofpacket
	);

	DE4_SOPC_addr_router_002 addr_router_002 (
		.sink_ready         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                            //          .valid
		.src_data           (addr_router_002_src_data),                                                             //          .data
		.src_channel        (addr_router_002_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                       //          .endofpacket
	);

	DE4_SOPC_addr_router_002 addr_router_003 (
		.sink_ready         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                             //          .valid
		.src_data           (addr_router_003_src_data),                                                              //          .data
		.src_channel        (addr_router_003_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                        //          .endofpacket
	);

	DE4_SOPC_addr_router_002 addr_router_004 (
		.sink_ready         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                            //          .valid
		.src_data           (addr_router_004_src_data),                                                             //          .data
		.src_channel        (addr_router_004_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                       //          .endofpacket
	);

	DE4_SOPC_addr_router_002 addr_router_005 (
		.sink_ready         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                             //          .valid
		.src_data           (addr_router_005_src_data),                                                              //          .data
		.src_channel        (addr_router_005_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                        //          .endofpacket
	);

	DE4_SOPC_addr_router_006 addr_router_006 (
		.sink_ready         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (addr_router_006_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_006_src_valid),                                                    //          .valid
		.src_data           (addr_router_006_src_data),                                                     //          .data
		.src_channel        (addr_router_006_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_006_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_006_src_endofpacket)                                               //          .endofpacket
	);

	DE4_SOPC_addr_router_006 addr_router_007 (
		.sink_ready         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_007_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_007_src_valid),                                                   //          .valid
		.src_data           (addr_router_007_src_data),                                                    //          .data
		.src_channel        (addr_router_007_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_007_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_007_src_endofpacket)                                              //          .endofpacket
	);

	DE4_SOPC_id_router id_router (
		.sink_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                              //       src.ready
		.src_valid          (id_router_src_valid),                                                              //          .valid
		.src_data           (id_router_src_data),                                                               //          .data
		.src_channel        (id_router_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                         //          .endofpacket
	);

	DE4_SOPC_id_router_001 id_router_001 (
		.sink_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                     //       src.ready
		.src_valid          (id_router_001_src_valid),                                                     //          .valid
		.src_data           (id_router_001_src_data),                                                      //          .data
		.src_channel        (id_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                //          .endofpacket
	);

	DE4_SOPC_id_router_002 id_router_002 (
		.sink_ready         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                  //       src.ready
		.src_valid          (id_router_002_src_valid),                                                  //          .valid
		.src_data           (id_router_002_src_data),                                                   //          .data
		.src_channel        (id_router_002_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                             //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_003 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_peripheral_clk),                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                        //       src.ready
		.src_valid          (id_router_003_src_valid),                                                        //          .valid
		.src_data           (id_router_003_src_data),                                                         //          .data
		.src_channel        (id_router_003_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                   //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_004 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                                //       src.ready
		.src_valid          (id_router_004_src_valid),                                                                //          .valid
		.src_data           (id_router_004_src_data),                                                                 //          .data
		.src_channel        (id_router_004_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                           //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_005 (
		.sink_ready         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_peripheral_clk),                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                      //       src.ready
		.src_valid          (id_router_005_src_valid),                                                      //          .valid
		.src_data           (id_router_005_src_data),                                                       //          .data
		.src_channel        (id_router_005_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                 //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_006 (
		.sink_ready         (sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sys_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_peripheral_clk),                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                 //       src.ready
		.src_valid          (id_router_006_src_valid),                                                 //          .valid
		.src_data           (id_router_006_src_data),                                                  //          .data
		.src_channel        (id_router_006_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                            //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_007 (
		.sink_ready         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                         //       src.ready
		.src_valid          (id_router_007_src_valid),                                                         //          .valid
		.src_data           (id_router_007_src_data),                                                          //          .data
		.src_channel        (id_router_007_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                    //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_008 (
		.sink_ready         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                 //       src.ready
		.src_valid          (id_router_008_src_valid),                                                 //          .valid
		.src_data           (id_router_008_src_data),                                                  //          .data
		.src_channel        (id_router_008_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                            //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_009 (
		.sink_ready         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                 //       src.ready
		.src_valid          (id_router_009_src_valid),                                                 //          .valid
		.src_data           (id_router_009_src_data),                                                  //          .data
		.src_channel        (id_router_009_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                            //          .endofpacket
	);

	DE4_SOPC_id_router_010 id_router_010 (
		.sink_ready         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                         //       src.ready
		.src_valid          (id_router_010_src_valid),                                                         //          .valid
		.src_data           (id_router_010_src_data),                                                          //          .data
		.src_channel        (id_router_010_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                    //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_011 (
		.sink_ready         (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (peripheral_clock_crossing_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sys_clk),                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                                 //       src.ready
		.src_valid          (id_router_011_src_valid),                                                                 //          .valid
		.src_data           (id_router_011_src_data),                                                                  //          .data
		.src_channel        (id_router_011_src_channel),                                                               //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                            //          .endofpacket
	);

	DE4_SOPC_id_router_003 id_router_012 (
		.sink_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (ext_clk),                                                                       //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                       //       src.ready
		.src_valid          (id_router_012_src_valid),                                                       //          .valid
		.src_data           (id_router_012_src_data),                                                        //          .data
		.src_channel        (id_router_012_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                  //          .endofpacket
	);

	DE4_SOPC_addr_router_008 addr_router_008 (
		.sink_ready         (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (peripheral_clock_crossing_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_peripheral_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_008_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_008_src_valid),                                                                //          .valid
		.src_data           (addr_router_008_src_data),                                                                 //          .data
		.src_channel        (addr_router_008_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_008_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_008_src_endofpacket)                                                           //          .endofpacket
	);

	DE4_SOPC_id_router_013 id_router_013 (
		.sink_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_peripheral_clk),                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                               //       src.ready
		.src_valid          (id_router_013_src_valid),                                               //          .valid
		.src_data           (id_router_013_src_data),                                                //          .data
		.src_channel        (id_router_013_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                          //          .endofpacket
	);

	DE4_SOPC_id_router_013 id_router_014 (
		.sink_ready         (sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sw_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_peripheral_clk),                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                              //       src.ready
		.src_valid          (id_router_014_src_valid),                                              //          .valid
		.src_data           (id_router_014_src_data),                                               //          .data
		.src_channel        (id_router_014_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                         //          .endofpacket
	);

	DE4_SOPC_id_router_013 id_router_015 (
		.sink_ready         (pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pb_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_peripheral_clk),                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                              //       src.ready
		.src_valid          (id_router_015_src_valid),                                              //          .valid
		.src_data           (id_router_015_src_data),                                               //          .data
		.src_channel        (id_router_015_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                         //          .endofpacket
	);

	DE4_SOPC_id_router_013 id_router_016 (
		.sink_ready         (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_peripheral_clk),                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                     //       src.ready
		.src_valid          (id_router_016_src_valid),                                                     //          .valid
		.src_data           (id_router_016_src_data),                                                      //          .data
		.src_channel        (id_router_016_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (5),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (13),
		.VALID_WIDTH               (13),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (pll_sys_clk),                    //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (80),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (13),
		.VALID_WIDTH               (13),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (pll_sys_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (13),
		.VALID_WIDTH               (13),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_002 (
		.clk                    (pll_sys_clk),                           //       clk.clk
		.reset                  (rst_controller_reset_out_reset),        // clk_reset.reset
		.cmd_sink_ready         (addr_router_002_src_ready),             //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_002_src_valid),             //          .valid
		.cmd_sink_data          (addr_router_002_src_data),              //          .data
		.cmd_sink_channel       (addr_router_002_src_channel),           //          .channel
		.cmd_sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.cmd_src_ready          (limiter_002_cmd_src_ready),             //   cmd_src.ready
		.cmd_src_data           (limiter_002_cmd_src_data),              //          .data
		.cmd_src_channel        (limiter_002_cmd_src_channel),           //          .channel
		.cmd_src_startofpacket  (limiter_002_cmd_src_startofpacket),     //          .startofpacket
		.cmd_src_endofpacket    (limiter_002_cmd_src_endofpacket),       //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_demux_010_src1_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_002_rsp_src_ready),             //   rsp_src.ready
		.rsp_src_valid          (limiter_002_rsp_src_valid),             //          .valid
		.rsp_src_data           (limiter_002_rsp_src_data),              //          .data
		.rsp_src_channel        (limiter_002_rsp_src_channel),           //          .channel
		.rsp_src_startofpacket  (limiter_002_rsp_src_startofpacket),     //          .startofpacket
		.rsp_src_endofpacket    (limiter_002_rsp_src_endofpacket),       //          .endofpacket
		.cmd_src_valid          (limiter_002_cmd_valid_data)             // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (13),
		.VALID_WIDTH               (13),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_003 (
		.clk                    (pll_sys_clk),                           //       clk.clk
		.reset                  (rst_controller_reset_out_reset),        // clk_reset.reset
		.cmd_sink_ready         (addr_router_004_src_ready),             //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_004_src_valid),             //          .valid
		.cmd_sink_data          (addr_router_004_src_data),              //          .data
		.cmd_sink_channel       (addr_router_004_src_channel),           //          .channel
		.cmd_sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.cmd_src_ready          (limiter_003_cmd_src_ready),             //   cmd_src.ready
		.cmd_src_data           (limiter_003_cmd_src_data),              //          .data
		.cmd_src_channel        (limiter_003_cmd_src_channel),           //          .channel
		.cmd_src_startofpacket  (limiter_003_cmd_src_startofpacket),     //          .startofpacket
		.cmd_src_endofpacket    (limiter_003_cmd_src_endofpacket),       //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_demux_010_src3_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_demux_010_src3_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_demux_010_src3_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_demux_010_src3_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_demux_010_src3_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_demux_010_src3_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_003_rsp_src_ready),             //   rsp_src.ready
		.rsp_src_valid          (limiter_003_rsp_src_valid),             //          .valid
		.rsp_src_data           (limiter_003_rsp_src_data),              //          .data
		.rsp_src_channel        (limiter_003_rsp_src_channel),           //          .channel
		.rsp_src_startofpacket  (limiter_003_rsp_src_startofpacket),     //          .startofpacket
		.rsp_src_endofpacket    (limiter_003_rsp_src_endofpacket),       //          .endofpacket
		.cmd_src_valid          (limiter_003_cmd_valid_data)             // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (84),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (13),
		.VALID_WIDTH               (13),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_004 (
		.clk                    (pll_sys_clk),                           //       clk.clk
		.reset                  (rst_controller_reset_out_reset),        // clk_reset.reset
		.cmd_sink_ready         (addr_router_007_src_ready),             //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_007_src_valid),             //          .valid
		.cmd_sink_data          (addr_router_007_src_data),              //          .data
		.cmd_sink_channel       (addr_router_007_src_channel),           //          .channel
		.cmd_sink_startofpacket (addr_router_007_src_startofpacket),     //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_007_src_endofpacket),       //          .endofpacket
		.cmd_src_ready          (limiter_004_cmd_src_ready),             //   cmd_src.ready
		.cmd_src_data           (limiter_004_cmd_src_data),              //          .data
		.cmd_src_channel        (limiter_004_cmd_src_channel),           //          .channel
		.cmd_src_startofpacket  (limiter_004_cmd_src_startofpacket),     //          .startofpacket
		.cmd_src_endofpacket    (limiter_004_cmd_src_endofpacket),       //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_demux_001_src3_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_demux_001_src3_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_demux_001_src3_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_demux_001_src3_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_004_rsp_src_ready),             //   rsp_src.ready
		.rsp_src_valid          (limiter_004_rsp_src_valid),             //          .valid
		.rsp_src_data           (limiter_004_rsp_src_data),              //          .data
		.rsp_src_channel        (limiter_004_rsp_src_channel),           //          .channel
		.rsp_src_startofpacket  (limiter_004_rsp_src_startofpacket),     //          .startofpacket
		.rsp_src_endofpacket    (limiter_004_rsp_src_endofpacket),       //          .endofpacket
		.cmd_src_valid          (limiter_004_cmd_valid_data)             // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (57),
		.PKT_DEST_ID_L             (56),
		.PKT_TRANS_POSTED          (43),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (59),
		.ST_CHANNEL_W              (4),
		.VALID_WIDTH               (4),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_005 (
		.clk                    (pll_peripheral_clk),                 //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_008_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_008_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_008_src_data),           //          .data
		.cmd_sink_channel       (addr_router_008_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_008_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_008_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_005_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_005_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_005_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_005_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_005_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_008_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_008_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_008_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_008_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_008_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_008_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_005_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_005_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_005_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_005_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_005_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_005_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_005_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (61),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (55),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURSTWRAP_H           (60),
		.PKT_BURSTWRAP_L           (58),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.ST_DATA_W                 (71),
		.ST_CHANNEL_W              (13),
		.OUT_BYTE_CNT_H            (56),
		.OUT_BURSTWRAP_H           (60),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (pll_sys_clk),                         //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_n),                          // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (pll_sys_clk),                       //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_in2  (1'b0),                              // (terminated)
		.reset_in3  (1'b0),                              // (terminated)
		.reset_in4  (1'b0),                              // (terminated)
		.reset_in5  (1'b0),                              // (terminated)
		.reset_in6  (1'b0),                              // (terminated)
		.reset_in7  (1'b0),                              // (terminated)
		.reset_in8  (1'b0),                              // (terminated)
		.reset_in9  (1'b0),                              // (terminated)
		.reset_in10 (1'b0),                              // (terminated)
		.reset_in11 (1'b0),                              // (terminated)
		.reset_in12 (1'b0),                              // (terminated)
		.reset_in13 (1'b0),                              // (terminated)
		.reset_in14 (1'b0),                              // (terminated)
		.reset_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk        (pll_peripheral_clk),                 //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.clk        (ext_clk),                            //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	DE4_SOPC_cmd_xbar_demux cmd_xbar_demux (
		.clk                (pll_sys_clk),                       //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)    //           .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (pll_sys_clk),                            //        clk.clk
		.reset               (rst_controller_reset_out_reset),         //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket)    //           .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (pll_sys_clk),                           //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_002_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_002_cmd_src_channel),           //           .channel
		.sink_data          (limiter_002_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_002_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_002_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_002_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //           .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_003 cmd_xbar_demux_003 (
		.clk                (pll_sys_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_002 cmd_xbar_demux_004 (
		.clk                (pll_sys_clk),                           //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_003_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_003_cmd_src_channel),           //           .channel
		.sink_data          (limiter_003_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_003_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_003_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_003_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //           .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_003 cmd_xbar_demux_005 (
		.clk                (pll_sys_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_005_src_ready),             //      sink.ready
		.sink_channel       (addr_router_005_src_channel),           //          .channel
		.sink_data          (addr_router_005_src_data),              //          .data
		.sink_startofpacket (addr_router_005_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_005_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_005_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_003 cmd_xbar_demux_006 (
		.clk                (pll_sys_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_006_src_ready),             //      sink.ready
		.sink_channel       (addr_router_006_src_channel),           //          .channel
		.sink_data          (addr_router_006_src_data),              //          .data
		.sink_startofpacket (addr_router_006_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_006_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_006_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_002 cmd_xbar_demux_007 (
		.clk                (pll_sys_clk),                           //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_004_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_004_cmd_src_channel),           //           .channel
		.sink_data          (limiter_004_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_004_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_004_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_004_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_007_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_007_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_007_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_007_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_007_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_007_src0_endofpacket)    //           .endofpacket
	);

	DE4_SOPC_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (pll_sys_clk),                           //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_mux_001 cmd_xbar_mux_001 (
		.clk                 (pll_sys_clk),                           //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_006_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_006_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_006_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_006_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_007_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_007_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_007_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_007_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (pll_sys_clk),                           //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_mux_010 cmd_xbar_mux_010 (
		.clk                 (pll_sys_clk),                            //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_010_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_010_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_010_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_010_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_010_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_010_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src10_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),    //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_003_src0_ready),          //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_003_src0_valid),          //          .valid
		.sink2_channel       (cmd_xbar_demux_003_src0_channel),        //          .channel
		.sink2_data          (cmd_xbar_demux_003_src0_data),           //          .data
		.sink2_startofpacket (cmd_xbar_demux_003_src0_startofpacket),  //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),    //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_004_src0_ready),          //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_004_src0_valid),          //          .valid
		.sink3_channel       (cmd_xbar_demux_004_src0_channel),        //          .channel
		.sink3_data          (cmd_xbar_demux_004_src0_data),           //          .data
		.sink3_startofpacket (cmd_xbar_demux_004_src0_startofpacket),  //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_004_src0_endofpacket),    //          .endofpacket
		.sink4_ready         (cmd_xbar_demux_005_src0_ready),          //     sink4.ready
		.sink4_valid         (cmd_xbar_demux_005_src0_valid),          //          .valid
		.sink4_channel       (cmd_xbar_demux_005_src0_channel),        //          .channel
		.sink4_data          (cmd_xbar_demux_005_src0_data),           //          .data
		.sink4_startofpacket (cmd_xbar_demux_005_src0_startofpacket),  //          .startofpacket
		.sink4_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)     //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux rsp_xbar_demux (
		.clk                (pll_sys_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (pll_sys_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (pll_sys_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (pll_peripheral_clk),                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_003 rsp_xbar_demux_004 (
		.clk                (pll_sys_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_003 rsp_xbar_demux_005 (
		.clk                (pll_peripheral_clk),                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_003 rsp_xbar_demux_006 (
		.clk                (pll_peripheral_clk),                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_003 rsp_xbar_demux_007 (
		.clk                (pll_sys_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_003 rsp_xbar_demux_008 (
		.clk                (pll_sys_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_003 rsp_xbar_demux_009 (
		.clk                (pll_sys_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux_010 rsp_xbar_demux_010 (
		.clk                (pll_sys_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_010_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_010_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_010_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_010_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_010_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_010_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_010_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_010_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_010_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_010_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_010_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_010_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_010_src3_endofpacket),   //          .endofpacket
		.src4_ready         (rsp_xbar_demux_010_src4_ready),         //      src4.ready
		.src4_valid         (rsp_xbar_demux_010_src4_valid),         //          .valid
		.src4_data          (rsp_xbar_demux_010_src4_data),          //          .data
		.src4_channel       (rsp_xbar_demux_010_src4_channel),       //          .channel
		.src4_startofpacket (rsp_xbar_demux_010_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (rsp_xbar_demux_010_src4_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_003 rsp_xbar_demux_011 (
		.clk                (pll_sys_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_003 rsp_xbar_demux_012 (
		.clk                (ext_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (pll_sys_clk),                           //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (pll_sys_clk),                           //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (crosser_004_out_ready),                 //     sink3.ready
		.sink3_valid          (crosser_004_out_valid),                 //          .valid
		.sink3_channel        (crosser_004_out_channel),               //          .channel
		.sink3_data           (crosser_004_out_data),                  //          .data
		.sink3_startofpacket  (crosser_004_out_startofpacket),         //          .startofpacket
		.sink3_endofpacket    (crosser_004_out_endofpacket),           //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (crosser_005_out_ready),                 //     sink5.ready
		.sink5_valid          (crosser_005_out_valid),                 //          .valid
		.sink5_channel        (crosser_005_out_channel),               //          .channel
		.sink5_data           (crosser_005_out_data),                  //          .data
		.sink5_startofpacket  (crosser_005_out_startofpacket),         //          .startofpacket
		.sink5_endofpacket    (crosser_005_out_endofpacket),           //          .endofpacket
		.sink6_ready          (crosser_006_out_ready),                 //     sink6.ready
		.sink6_valid          (crosser_006_out_valid),                 //          .valid
		.sink6_channel        (crosser_006_out_channel),               //          .channel
		.sink6_data           (crosser_006_out_data),                  //          .data
		.sink6_startofpacket  (crosser_006_out_startofpacket),         //          .startofpacket
		.sink6_endofpacket    (crosser_006_out_endofpacket),           //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (crosser_007_out_ready),                 //    sink12.ready
		.sink12_valid         (crosser_007_out_valid),                 //          .valid
		.sink12_channel       (crosser_007_out_channel),               //          .channel
		.sink12_data          (crosser_007_out_data),                  //          .data
		.sink12_startofpacket (crosser_007_out_startofpacket),         //          .startofpacket
		.sink12_endofpacket   (crosser_007_out_endofpacket)            //          .endofpacket
	);

	DE4_SOPC_cmd_xbar_demux_008 cmd_xbar_demux_008 (
		.clk                (pll_peripheral_clk),                    //        clk.clk
		.reset              (rst_controller_001_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_005_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_005_cmd_src_channel),           //           .channel
		.sink_data          (limiter_005_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_005_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_005_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_005_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_008_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_008_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_008_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_008_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_008_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_008_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_008_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_008_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_008_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_008_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_008_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_008_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_008_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_008_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_008_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_008_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_008_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_008_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_008_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_008_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_008_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_008_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_008_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_008_src3_endofpacket)    //           .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux_013 rsp_xbar_demux_013 (
		.clk                (pll_peripheral_clk),                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux_013 rsp_xbar_demux_014 (
		.clk                (pll_peripheral_clk),                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux_013 rsp_xbar_demux_015 (
		.clk                (pll_peripheral_clk),                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_demux_013 rsp_xbar_demux_016 (
		.clk                (pll_peripheral_clk),                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	DE4_SOPC_rsp_xbar_mux_008 rsp_xbar_mux_008 (
		.clk                 (pll_peripheral_clk),                    //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_008_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_008_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_008_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_013_src0_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_014_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_015_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_016_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (57),
		.OUT_PKT_BYTE_CNT_L            (55),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_ST_DATA_W                 (71),
		.ST_CHANNEL_W                  (13),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk               (pll_sys_clk),                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),     // clk_reset.reset
		.in_valid          (cmd_xbar_mux_002_src_valid),         //      sink.valid
		.in_channel        (cmd_xbar_mux_002_src_channel),       //          .channel
		.in_startofpacket  (cmd_xbar_mux_002_src_startofpacket), //          .startofpacket
		.in_endofpacket    (cmd_xbar_mux_002_src_endofpacket),   //          .endofpacket
		.in_ready          (cmd_xbar_mux_002_src_ready),         //          .ready
		.in_data           (cmd_xbar_mux_002_src_data),          //          .data
		.out_endofpacket   (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data          (width_adapter_src_data),             //          .data
		.out_channel       (width_adapter_src_channel),          //          .channel
		.out_valid         (width_adapter_src_valid),            //          .valid
		.out_ready         (width_adapter_src_ready),            //          .ready
		.out_startofpacket (width_adapter_src_startofpacket)     //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (57),
		.IN_PKT_BYTE_CNT_L             (55),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (60),
		.IN_PKT_BURSTWRAP_L            (58),
		.IN_ST_DATA_W                  (71),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (13),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk               (pll_sys_clk),                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid          (id_router_002_src_valid),             //      sink.valid
		.in_channel        (id_router_002_src_channel),           //          .channel
		.in_startofpacket  (id_router_002_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_002_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_002_src_ready),             //          .ready
		.in_data           (id_router_002_src_data),              //          .data
		.out_endofpacket   (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_001_src_data),          //          .data
		.out_channel       (width_adapter_001_src_channel),       //          .channel
		.out_valid         (width_adapter_001_src_valid),         //          .valid
		.out_ready         (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket (width_adapter_001_src_startofpacket)  //          .startofpacket
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (89),
		.BITS_PER_SYMBOL     (89),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (13),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (pll_sys_clk),                           //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (pll_peripheral_clk),                    //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src3_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src3_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src3_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src3_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src3_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (89),
		.BITS_PER_SYMBOL     (89),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (13),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (pll_sys_clk),                           //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (pll_peripheral_clk),                    //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src5_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src5_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src5_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src5_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src5_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (89),
		.BITS_PER_SYMBOL     (89),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (13),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (pll_sys_clk),                           //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (pll_peripheral_clk),                    //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src6_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src6_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src6_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src6_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src6_data),          //              .data
		.out_ready         (crosser_002_out_ready),                 //           out.ready
		.out_valid         (crosser_002_out_valid),                 //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_002_out_channel),               //              .channel
		.out_data          (crosser_002_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (89),
		.BITS_PER_SYMBOL     (89),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (13),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (pll_sys_clk),                            //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (ext_clk),                                //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src12_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src12_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src12_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src12_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src12_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src12_data),          //              .data
		.out_ready         (crosser_003_out_ready),                  //           out.ready
		.out_valid         (crosser_003_out_valid),                  //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_003_out_channel),                //              .channel
		.out_data          (crosser_003_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (89),
		.BITS_PER_SYMBOL     (89),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (13),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (pll_peripheral_clk),                    //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_sys_clk),                           //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_003_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_003_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_003_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_003_src0_data),          //              .data
		.out_ready         (crosser_004_out_ready),                 //           out.ready
		.out_valid         (crosser_004_out_valid),                 //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_004_out_channel),               //              .channel
		.out_data          (crosser_004_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (89),
		.BITS_PER_SYMBOL     (89),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (13),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (pll_peripheral_clk),                    //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_sys_clk),                           //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_005_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_005_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_005_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_005_src0_data),          //              .data
		.out_ready         (crosser_005_out_ready),                 //           out.ready
		.out_valid         (crosser_005_out_valid),                 //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_005_out_channel),               //              .channel
		.out_data          (crosser_005_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (89),
		.BITS_PER_SYMBOL     (89),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (13),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_006 (
		.in_clk            (pll_peripheral_clk),                    //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_sys_clk),                           //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_006_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_006_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_006_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_006_src0_data),          //              .data
		.out_ready         (crosser_006_out_ready),                 //           out.ready
		.out_valid         (crosser_006_out_valid),                 //              .valid
		.out_startofpacket (crosser_006_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_006_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_006_out_channel),               //              .channel
		.out_data          (crosser_006_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (89),
		.BITS_PER_SYMBOL     (89),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (13),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_007 (
		.in_clk            (ext_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_sys_clk),                           //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_012_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_012_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_012_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_012_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_012_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_012_src0_data),          //              .data
		.out_ready         (crosser_007_out_ready),                 //           out.ready
		.out_valid         (crosser_007_out_valid),                 //              .valid
		.out_startofpacket (crosser_007_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_007_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_007_out_channel),               //              .channel
		.out_data          (crosser_007_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	DE4_SOPC_irq_mapper irq_mapper (
		.clk           (pll_sys_clk),                    //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_peripheral_clk),                 //       receiver_clk.clk
		.sender_clk     (pll_sys_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (pll_peripheral_clk),                 //       receiver_clk.clk
		.sender_clk     (pll_sys_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

endmodule
