package rmap_target_write_command_data_data_pkg is
	
end package rmap_target_write_command_data_data_pkg;

package body rmap_target_write_command_data_data_pkg is
	
end package body rmap_target_write_command_data_data_pkg;
