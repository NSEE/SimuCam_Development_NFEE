library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity comm_spw_codec_extenal_loopback_ent is
	port(
		clk_i : in std_logic;
		rst_i : in std_logic
	);
end entity comm_spw_codec_extenal_loopback_ent;

architecture RTL of comm_spw_codec_extenal_loopback_ent is
	
begin

end architecture RTL;
