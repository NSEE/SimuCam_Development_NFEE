// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:54:03 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CDXFU6jVfoh9snNx9zfFjbRKroK2D7HsNkd1liSUVwzCyB+XNaTtu6e0yOE9iRNU
qppMwj4XpUqd1G+TLnMr+3CY8alEbppnb8bY/MUCH4l36CwW5DeR5hjbLmkc03Nf
fKwzOj/U6dEGmSnrDdMdYUgjxcl3Ck/CZZjZ9oiEBNU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17008)
NBkaDv9aDH8QQzFaYXyUiEMxf9hsTAZfNk6g0LVNrOIhyNPXhegDgD2ZGMz8leoU
F9eTV6wgpHiKzJ6ZMTxex9szunb4dCraHRojYv2nokpx/9thyVwDc/CL8w1Ea7qH
phfQrWjy6F19vt0FjZgTyuLqIB/D3JRLXZHFKKsV7XNq0luWsKQ5pg4U+6sfUI3S
nweLc6BQjs11An8wrTH8JFfaLO0uiYdp1STP8C8tZ6TuJujbE9JVbL2OonlUrFXX
D3B2qI7dDqpOgDRNGszozii88r+/ewCliDculkqkfgO0WXrx8G20pf9MfqsA6LzB
VY/vmWfVNTn/SclzgndtvgGk0MqFeQZLvyfNESwOPmKK2ydD0N7w0cBSAVJf2SXf
ZCCWN2kCUOlr22GXgBw/YnmMBcX0xarTTRN86WwtmYbi57UigBIz3culvEVjnDB3
ZBw1OZMvS3+uNijW5FzDfDnPfgZ9FZpbgklZBjcmRhC2ukBMg8694wRmuyXpA1B1
4uw7ldbire66me38eSqXIP6Nr2Rt2aQIgWkN53h2imXZvU09mFc/IMTonc09zIUY
7cSm1Xu3S5qHoRqaj//0xUI0LXrbO1VW2eVDJHgAsVWfOLR2CG5G7nuVKn6+Ejqx
HKLN8KwW6X3SR3/Bf6Nf3dtec4ZBin8E1pSmZ9PTIR7rAKzR0XbcC8P22woL1p5M
MuffZC+WRuOrFk/3fdPqlzmPxCmTZBTJt5F9jhLzYWjcgkFVq+G3hCI/czpYBnDo
YgSNsYPLuv+eSdIuKQpIzF6JYJDajJCQO6ewfAaEleikpTVDy7wHJtL5oTSuZDrz
9FUOHG+Hws5K+8hbO4HkHVCjgiEg31VCVO2f8bmH2ghwfgEi72aFXKygmk/gHFtf
h9opZgGeI4iyXDjgq9pbdA+/atuGuyFlmiorywuSIUixhJqhJ3ECyMeA+zbBvref
+efCHcmgdDF3o5jLM0k5TlHpIbOETqfQ3djHgcI7SuGs/QMUnl5ky6Q7R0/f4/qg
VRIF5iBUWCnr8xcP4y1wU8Qo8FQS48n2kd1BvnK4bWsjWJkm5LSeA5ZtKSEeIGoN
r2bh1nbN+ZQgF0w5mLUTA76Tyl0Hx4qh1gFRsrIGilZwj/shxCffJ8GPssaLTbAX
NB/0gjpj6s0dINT3UtX7NK3pYcFkw60OpQmCAq+PExUA/VvLqd9Jsd6TKvj7S0Ee
e0jNBNRqQhuczo32DVcpRewYhTLqKUiupPp5N09l6/BEL/CAlqfkY6Eul0aQMhEj
yToLYtOCdSWPhQHo7EJ5SevlL4Xma5cYomhbVk71iCQegRQpL5MchxkywEMrqcw7
7xDcHc7wcwhMkajoFChQqaF9AjQrY9KkfoYfWvs5uoggeN3Cm/m5CclC6xCuPBXY
xWg3CTt0kcBeU4AzEh1+1aMobm9r5EgyjwActH5wMSQhn02zhU43Ar2XTBqJ8I3S
BRTeOrafwcqaePKVxufV5wgtKPlH9xdV7zT7nmKOplVDDKxViCbZhrgD2QShrlr9
Xvz0Yso7R6ta8QVTXdOXX0Ni1nSbdiugQl46Fx5qOmRvnG9Jag+jcV58A3Pl80+V
MBBU3ldAcDb2NV6TN+9ovQLT+vmOBJ6YreiLiAZnOMJ3k0a098/+TjZyxv6D8ppp
P5OidTPydv02Bfp91fqe3P5X8ZgGAX53vXJQO4tsbPcqH6z03HY9TavYQ9faqmN5
oKLJk/hKQdhD30+z3TmB9FG26wQMt7xLKMzvsrh/V0vmuIabcadjKWiVpS76UuxY
UNJX+KK1WF/DWlOhJNrcy8xVtxgvF1riOe5LoylyRfQ8THfVjv4s6p+X98rmmzrz
tyX2ek4yY2e9Qf7qyItp+gzIum39i/9jxlSWQ22lZ+c/vHNzGyUPQ6df2YLQ7ar0
FuwSGcOSKKum9o5Sdnf7B1T9RYhvTzrwJRhRhvPOgXv5bKDiDE0MsIMWU/QpEafs
YhBoaZqytbqwTBy5YjMC8ypEwTbeus8KPtZX4mdbDnG7+4JNLYUz5KN9cWSAVTGC
xXqU84ttNVpjGhcJ97gSrapGjaq4drnmFPbX4t96batgH8MXGv80JX8X4vyzsqE3
UsqjsExs5Ti+8T0XjFkzO+kAZV76iRoD+GSIDmlzTxEdqaVP5Vu3QhjoavRjXGn9
v7yx4PzIp8yYDNV4yFBLgwxy6joGw5IFQgzGTlqDx19vl5qXRHkUPDydHV4NwlrR
gRqx4EBXytp07mSDKXx9QeudyxtkjCOLbTB7ZoAVhP3mWgv3uy06JlGHqaKJkys6
u/5F2TDLYzUO0MrMbF1VCDecet4gNKNhqH+njPKQb0+jgodTLEB4fCD/C7A2dYsY
Fhrs79L/550Rd9+MAAffk3l9jjmf1mRWzkHzgb3Ct9vn4Z0awSVUSVak89ejRJOc
Ex89BSWPa/BWhz7XrPVggpfB33l7cXPslD7fexhwmeQmsJ8ixEEvx+dHE7thjCaH
l6totzGHHwrM9qcAsfZ/Wa+JlPkJB+e5LvYX1UAmJGFP55eIcsr1Lf59WRfCAqEF
ulV8UrYnmKLV4b7iuiTGPJKF9B50bc/asUGGp9I/6wR+KtPnN8WwQtrACXUiX+N6
cSscerkZWjDKPa/83IU4GyDNr+Qcp+fXcOW2DIAzaUHcdu0q6lfoBZ/A+jTce3TQ
OKm5cH3DcG7hzd08ZAFCR+Y9W0UEj9RERCc22yyisO8cJp/amzTnFvJPfvnml4DM
XocCnVs7MclM7+pp1uqUeywW14XJANsOieFii/3sgn0gRusJe4XIoU363tRq6jgm
pJTBjEg2jAClg6hkU9ru2+6i3KhHEVGy1BjXpUqQq0stnlnuRJkSqOSglGnRIlro
s7EblJHxgBjgsGpPJPe92gvCs4ZEEszbuJp9F2AtpPWd7fRIy2P02Nh6ZTqTfUkA
V/8sp3ry9O4Ov2fsCSD+AxhYCmPPsoL3YkHhLYijf0dlrGOUl+WcfiRI0gYUMVu1
y56MbXPIfe10UNHpswlJ1aNExPiGrd3gcMDkIHTH1Ox8FrnM0f/T5qhsBhQa0HSF
3Fuk48SneY8CYyT8tKdr8J6/Xjp/pIiGmvdIEkvxm/zXoAfLA8g9mu9HZlkmvyfU
JuwS7Abkc3dg/P+6GxHzO5tcDPIsT1T8ltVkqZf6czx1GUlw6uB9o9gugw7c87cW
eUjgWGmNSAgsof/KG5mfblSUBWQn1x8b9x41PzRruajaOu/OeJETJipEjp2w9Cgq
5rXQPk9FEt2NweOPcUyfOsP78hFXcsigJcj1stcCojWcXNIgeYiZSkb88ct66liQ
efF2KASX0uMi1CJNidqnvel9W96fQlPqkHFo9JtrrLOrEtqN148q8nCGD9+1DnM+
C9IBp+VkznwtY3FhXuKbVVFEfOLbJvlW8YGO/BLyIIRvIij0ysufen9srfq5F6zg
tzdrDz+N+OYRukdPgloGxW1AhohJz/1itASAM9jWqbuKqmSMutqIdRHWD+FMBEZB
sktxj2HP8aUxVuZbgIE8ugdYIBWMgz6yoS5sLq2SblfI/+lqKxPJ0I1USAIy3RJy
3oCNLwG3WJ+z2Rhjwz6uIL/gx+uVrsPojlW8BFITD1xMWN2ELgBW+ZzTIW023By8
0JLfuA/c2uDMwa+16rZ5vKpu5n6Tbx8yzh+EPo+Ypmb2brx6lr3mu0I3lXszYBuX
XqfXwHOqquiA0J6oTxfpuA/vWNLjtSy905Ns9ek+q4eYEIkd9jGbyu627l42qQGm
lmJ45z1nZCkUmR/dWXgbnOAn2O5WEmMayVYDNoL7FJfncOIIXc+hPK87gq/Rxt01
7Yx6Gn1FVdaDXL9/T1fZl2LEMqEUHuehk7Zmyge0ONgOgPdFkUlN5P/ls/NzlDs1
kICQNKyymup+V3GAXBZ9HcjVEWRQcL2Zw+5gBnZPdkWY8gRU2MNVK4cUDfMFh6cN
AZvZtInz+lMm0QhV7uO6jaUJoV5PegLLqKGQZ63OY+LxLiLU8ZqHZ159tlyGq433
tpNrcRyTxJrXlah2v+WbGLpj9RykORF4GMfosxWsPdqf6owbSty13YGUUwZVShsT
X2GKD90fLlut4ivFsiNBRPqKO6eyzG75RGJZ7vSNmYkN77kJf6lmJz4i07S9SiaF
loJrvDL+TPHeb7HowjslPSkMrLp5Flxyw603xysP9971VPl8FI/YEiRMeIT0KYn5
b+2aPJc8CDo3unkmH8nb/JIimp5usnfYEivbCzS33G3XcDLFPT7play5TiKTuBDz
KlkI7n92y+iWliPOl6jBHqnV2Y6u8yr6pIQigy/iXoSfSTxhCfncQmfSqZ4PmA1F
k1Y/bieuR7xH4uVctwSU9aZ6t+l38eP4v97dRmJYDGAzcygo/1EpwPvP3nM4Yv5T
Y01F9rSDQDf/HTgxYjrkxq3kSn3yVyn8UgkdePDzYxv7hjS0xCsskQ4GjVSSGV3j
/teSh7+D7G+DE7fPtp1NVPS/tSJqibtxwugYwILUPl+gIuIUcqsZujS47vRAm3zj
jFRXdhQHulUlVcW5UCED6xoeyAykYzFmdiytpCm5SjuFzK7likKZzQnGKQvbjt59
GsTW0knnOCo498pZ0YovcNn1YS8B0pmTUQsVQZ7aAloVuEVEPZ9ddqK3TZpM6FJj
cbMNpzS9aYOF/Rnsdr8ZTt27gT+ACFX3H7+Itrn6L4uB7sNA4RL2Fq00EPVo5DW1
VrE1tUkbWK5I/F7Zn6btGKMgMtauyNrPnevt20r0uqyIuh9z04gCoyUt0u0IgYA+
by2FV6vF6CKeGGLps8Gzgfmoj2ZJZd4DEAjyRLLyFWwrhd6lh1XnC2D9SwJ6jsxh
0ieKjopoXgt0vTqxVtGxUwwkwuCqQrczQKLW6+BXnm0ftXD/iBj5NvtsS7s2/8iN
x5fZOydc9v181MGHooT4m/zdv65k7nfJzOgJ+GRoaxAIEOt6R5xYGFfmF90dNTZf
3mh7+WR5TX8S9GFTVrK+U7EcPSfJnCHlVj4zpi7sZGO+ZE0z6KKCxW2kIe46+Jiu
TejBJH/oC6B+zkQaCzJcqRXfHuBAj8EFOBo1e8NJoD4+gGp3JfTqhSVY+B/J8Umo
/LUsepmODW5p53rvmJKNAXkZbKhVxOQpzrI0nAI4hnffrW5ItnoAlxb2WGw/lZr/
jWh7SaQ0HHbHSwIXM/omEq9PmcnQBaOMPhNjaEqEMe1hIrfnq6doSBvAq9p58N6v
yiaarKiHoEEIztI7hakBZmxqSLOTcOpKu3xfNz3gX3Z7Xcn0MFTVbl2owaDEldqn
eU42MVQ9LQmvltnX85wiYqZXOMawblNVwZWnw5z41cbDJVy+ZkBSTTdk4Vyk8nE1
ATLhtWJlTHML1woR0Xl+hFp7jDKGsXSVOfQHkcG3mrFcIGCoKeTDvp2wgA0UN4ZB
MVZR7ffnKpP+FEdD1Ws8No+Kn0KhGX2de6OyJoPHhCUtyKkANA1bm9aE3QM3VJB5
Dwe9V7QgqJT9qzSV7RnnYb8KvVOcffNeL5gY1N91azkL5wl9NnFwqMzHyPe0DUPt
gVETmIREgLRU5UZwRZXyaMBVkn63mjS49QVxChlBZolqnh086blA8YQFaUm3sE1k
fHQZs2uOi5LQWr2BE3tdeD5U1MdDGCIx6jICA30EaYsTdRgu+KzLUeM5R2fMUShL
/HV9k7Wf5rY9Bp0LHuJp8ssG9txhf1z9rHJYqbOEuMKd9CxNPx3U/Exj0Mgnx/5q
fSjAg6cssHy8PoAjLy5mWwy+pNotlh+WMOsS+lE9WwFwLtNu4d4495nY42ItOorP
XXy5ca7NUKTkAG+gwKxgSwXuW/LhmTsenBWifTS4WWPGrceRUmjoWlsLfw+VJEwX
PtGNncgxPZqivCgRiMRwxN+us6hgCmDNw04o84dgj6dUnqPNsDIGmkeFXJws9muL
/inVaw3NArx6wkkGEbVFNY13wrvDEQoAQHsNWV7v+UNXJ2yV0mDdTAvyrzlDTtPZ
xUo66VIuIdLTS6iZwxg3UZI4wLQj5kglTOtfW26OJk58somAS6FcXev+0dZd/5El
Z6zj3Ax9+aSSgvqJeiQ3NTt1785xqrtKDhBnx5uLYWt0jhbOFpthAp/cUSq/lYYa
iYnt0Wan7z1dXh6zYtrra8to3MdIdl3DGPyyw/3q8DPC+4YctT3DwJiHJT8pUADr
zt7vTlhOn81ez9kdEL2IWZUi/JjyEtLyBu2cQ7N81t5/5Uc0LKwqpX/4f9+/Z7jj
g9relaqy7yYk5CzSz97NnDJN9tOZ6HYYICCDysxugSltcEbj4jIbegXQA1B6e0V9
H54C3dkZBk3UlR16S52z8KrJDkx3TyAX3i3RbvGXWJHv7RLyGxUE7jd35yZvqTX9
YkQ7Sqn131++k6LvGeg30GWWqknOQhaupCGtnF13qit+kc4e055yt8Apbx10dkF8
/Rek9yEfsh0c11ZMuS4ricUv8Qgwf00BX6WWuNA/E2p/ADJfAxkvVGwYd8cr4XmK
MtLEWX92tqhZ1tkuGze24aB3oskMBvhltcUqSh2CrjVHAJJQXJNIuYevWnq+yllY
4cOiJg+r5c7LHcK6gHJUmIYX15a+s29K35C3LUG3b08kvczj7sfrKOkWSNryzN8J
6UxKK3O34496jLhIk+nNJ88RFGDGozNNU2mNdk2/Ontz1EfyIzEGURP1pOPTuVoB
Y2O+FBp1tTzLBVdzTIJfBZWFlMFSriRJxgQwZINA8XSGZkiKyJNTTKfe26sFX/VS
a52tVBPtMbwxfc/fcdgo/yAf3Lzhe69z1vUg2ZhegUXWrMozo7mEBWEsowe5xuDH
4AlXjXXZ0xKjvslw09J+Cl3AaTtsBBl6YwJu0+Q7pUOBeJI/LrZZALeG4x/cE5xf
zzEYAC2ouUdPUiG7oh6/ySmMgQvNKljvmHtYid6FTQe291kERhKPkpj2kCh7XrVe
XOQhyW+ZEFI3RL4zpVNZmwfE6RqJlNX33JNEs6L/n+wtjXzFz9Fgd9lQg51ndNfe
2NlgWdP1vh8PmkfyTF7FcZniQwp8vvWGRDM7zB+4rrHAv8z8287y3JdubWHRU6QV
zVEyyKwmjL0pgXQwkyNKTIF0jIlGQoJD1o/hIZxQxFZp4kw3YNQ63x35iKXVcnKI
MnWjs6t7yG3ZTirCRUTlN6vpzIBjlHGBQUonnbDSG0JLKpKoGAY7jcy/wyIysQUk
k6PIdz0P7fm491cUGV4VhXkjAgnIUTDt1oMXdAol8dOwRj8aDvZBcs4gntVb2jiA
lJPFKxcvXm8jR13AHljc5+OL+mpZq+TinQIFcNdUxaf1FbwwVIpxJx40DluFotWu
HpplJrkRetePiuYkR36Ne5HJSIH11rzCK7O3Ed2l7W8eiQvwQYezfM0V8TwYCaB+
LmzhZYKygxAAM8XWdpnb8dqKh3szUsxvddelql/9zOXjG33rIpMSiMedly4nDMRG
ZiuAwTohfloshjc7zKs18ndxOa+eESeH3SEgEbvgFFhw8F2w+kl66Q7q7w7sU64q
PLH3J7cRMZFs0VSxo/fQB420KxQlMbz+OE7AA5UfCUUbDUCTCuMhdhZ00q+G4GrG
s0IELMGHFtTdWeszOLubdP5K41hBKy+MaKqUyjeuHoqGRyjobBw9xlXQvySH4Nbt
V/Z/3jcvBJ/8x1cyXZu3TtGimYqHdWPZ6jwJG1yiE8nBdMkWgV3T9eC9juIsvhpT
aUtszLr9jrZ65TWu1pepcSNsAVyXchGUif2kPX+rND8w9kk3Jxo+luULOor2/J5G
/Muy7SxKR7BTQUJh6vV8w4bZc3oxr7R0x4ZdA7EUJ1X0DWjDLigxCVbBpxNEwNjg
qjFp+NLUX1C4JbnEVAN4W93lZj7Sa0KUax+roICle36SLgWo39ovBSVrLh/f489M
CNbW0KP2a2TcvahZfSv6Cbh8SpQZLbLfvwqrLpuoFP9KvYM5ck8TsjwIynE8zCIy
bBcMMExlFP2Bywgxw6UlxtUCe9uU3V3zf2a3+QA4xo6mDHRmRYJGUZ3yHwlGmM7o
HX+EdI3GC8E8QqpDVlODdDN1vJAtnM9h8X8W1LXF6xi0ESRFg+EXWBypwmq5ABdt
tbANr8aC4T7jNIvHbMfuRnl2U1kx8kaaFuo4uoB74fypQ9sCNWQ9KdvBU22KssmZ
EjSCOurrsq1e5lrxubsekAYu+hbQf+dw7ysD5FcTiLZhBfVxRFd53bVUcmX0mvA6
QBQOkjzJ0aXl6sdT3Cr53W2nIcZm3j/t0BkHRWk0CR8JJEQLpuU+etu0Wilexz19
/nBtn0iJaiAMpr+56EFQMelXhAMLIk3lq412lI6jF6mnbsqChLvPrnceY0WDtqyl
T827ZPVQoSSzoSKp2CdMAkhhr1V2GqtkiMrjv5qQ8tL5qFC9uCnblCdyMg7iX0kK
PsIWr7XHprrYXQZK1nRmyU9xRZ1Ma0OeCrpoZOzBA185QCPcWWtQgkW6fkLimwy2
l2glvqi9hjcjLN9S54AeVXqlaf6L56Ayhknr/FW8N5P81l4nkdn/8MVfyTIfRai/
u2XbbRrGWoyxZUxDzCm8BcfN9EK5BIT51Nli93ViKcARPxikZ2K5H114jh5ipaWv
13BpnQDEnSFNlakeL8gwnB+3ve/FBO2N1nnp/TIjsJaB6PU2nhOw5cBylLUrHp2F
yCDIhWyApHyv34ncdAtZ9RbDNErwFRogdhOIiklG+w2wZOl/Y5xPu+4Ysq6+ERoy
iBrj85UVBYAoGDCGtF8ZkF/+JfwuM+rrgd/MoBe9r+h/vclMZ9KP01nyi2k8e1vl
5EXCgt3ZK1Ot5CX277vIvOA7X6Rs55JJVb+lgPWpchXZTeO+e36AQd8ZZf3JaIbd
2ytzuOvcIDlBwhkkEoxq02lq1z46AnZu2x6qdv1mRxbzaQjyWFVwzGt047NPoGAL
RgL5KspAbtkyaBV8hqe0/Lj8DLrs9O8pxjXi7wmchHW6uVaKcVN3bDDFtzByf6wE
93aE0BmAKipMBEaAZpdh60b9W+VbNAogCBfyPq7YzrKkiUGY0A9HOX1p9YiE0uNF
prm/7YsA0htxIDILbF2kEzYUe4KIaMb2yd/38DGNVffi6e0FnU4l9f4bgtHZ/5v7
Lxe/74UIPAVuteU4Og3pR9o7zc9tdMaiWcfmUXrSi1uLeHtdJTWR5JUjL/Ro3grX
YoE76U0QlXMW4MODx9bTmi6jWzhZd//frhcOKt9vpHlHi0gWdpOkO5j+5nLGbmxm
ZIoMXTfpUbkLBZwdxu1rtJMp5DaUEJUIMl+iQIur3Zc4jobvkeuDdoJHazrTJD8/
+xhPH1lONbcygtZ1elDAwGkHZrqIvZOJXqFrmcSLvYTHsKpHE3N1rNcbq6/7L4gp
3Mi8slH0sWk6raB9yGFSSHFuTDOMgO21blIGj5wvav3SOT/xcA0kx/47DGfbjdXi
Nu3MUqv4lQASWnaUfmFkWrfSfV3zyNxqEunCWZ0//0i8mSlWVIqO9UC5n/ZhPYdH
oKWOqxdLKiISSbv1mPUgfpTLSqG3Kqy544x5v6P5WAhM+7625+XdhwaJCKCpxTyN
V9ptNN3G4UWasuLkDnv+u5SP3qKGCNIay9IpDmSdIJzOxGpsoBNr2ZoSl3c1S1vt
7NXd4liVz2BaAUJ8/qNkYmfTJPdXRpQhlioC31TpA/lSAynDeOYmC6Q2y1GNPn0P
H6oueSp7vnGcutTMa0rhxNGJApCWHVtOHoVRzEmHltR+P5tXDZ61DEaOCwgcqJz0
fjLbuwzMgpYmP3R5dO+o1fGp88M9AUB0NjsdC60uhPEvBXmWSJG7i1JwVTuvXi/z
sOqYI712E1F8rw1vX2lgrmvOSE2pMlHLlswfsrjsRL1ltvibApXJznDaYniFYuX+
RC8bYjzGyl3u3uIwFzZN5BAkjTn9mAgo6FYy8RhEoqrDThAI8aNYzrM4G7crnmW/
nHV7NczL+Yww6fgRSBK2hxA+QLPIbvmegtj+NBeXsEWQ7HCRvL1WR3xQiSlWqFBg
Edu+udtpx+PstJP9zT1BVgBUcxzK9ocqI2L6JBgDvzXCq/VabPQ3Ukb4gHFOe0GT
CtaDx96xkg7sT+GeM1RTZvFRleClt/j0OopVv+UHx8mF+cAj8idyP2CutTi92DHZ
mp0XMOJiydBwnFhAYkfrHMS4a477siE8cOAafqbp8C9p3VpZPSP1lID558FF/djO
moXLP+g908NUK5qu01GAetS+m11ohYxSVZ6zI4tEIrNnZndH7qDgqRfGdQZ2J4Ku
XVVHaKVdUaJIg8azLw8m9pvtm35GFEAAddjoD2cJB+X5I4CQPE6H0gQ8l6KYrXl1
UV6srQ9jqs98UHXVQAKoGV08da/f6kXqesDQbpaYrVKTsBsHnLmCHqIzlzzAl24E
ZpWFmD7j0yViYXWxGhQx+FREQ3/zMFU+I8zpXgu6PRZVoFEpXI7zZlL/lQbsZu6/
1ch614kG0xDwNv0j5hBLuC3SDCBEanwyyy7gQAQbWFxjlxGhHmxQY8WnZIwgRrG8
qm3goq7l8a6til5L218utndrz/TrxAgbJrfmv42OYrFDQlCyxIFG1dHX1EMyLW2i
ZfSKw88uJQOZwr0tpK9HxPfEo2P4txYZ6/8hqpcWAvihO9q9kl3p1ZxbbO+/WJE8
6VQzxo3KIeXyjwIsHm1/CxZqFhMfzuGKgzZH/cv8JwKr/1wkk9o3LG2caW2Dimu7
YdmDnxAH3daWXhdw5FLyDFpF6W76Fuf0dMW6f1Wt+CZAuwH5ZmQa/dLCtMXmq2Bp
6Z6RUOc1pWu8noFxevNLpD+dB3TmVk9P+4gBuI+JIscVooG/xEX6IIeoQtD/qDh2
y0c9wEPA/MCw1rmAXmt5hzJT/Y1E0sAVVCXxw583JhsgzOnrnpnpKrw3zGdMf9LZ
6WRGr2Uoqee22f9U9cjxsURe5TD08IQg22gmaekp949/TVlpBNUfHjoSU9klSdxz
PAZ7+w3bzvew8Bja5Vf1Sv0nXatFC/Hbt/ZETP0ewbdNLswzBEBFjcBXB5yN8jDj
eH5/sKfS78rH6FCJBlq8bD+6rWIh+t4pq2mBdIdgciQEEe4hih6Bo0pKfHUNSqD/
/Z8fn17xYIq8LNUDC4qvB9kcfa48hyLVB/rQ6xuXML4VUw1YFVwQiAG0LVgvQ/PK
Vuvr++GsNsT5Gwoe0YMFSFLCCCH/ngxu2yu9wOf2ezxjuQIXT2pK+R6BeqglyJeQ
sW6OOxlfiEVF+iRF0FBslAppwR/IAxufRikn8s/nwE0VbaE4FkzSGFK3K0mpYC7H
jDfBYCrUaIvBxvdQdBhqzcdLtNCrKftz2eg2utNrXHHieuT0P/hMIzZSJqJ9mXHI
cLPOOlnwCr1KT9AhWrVO0kwb6LxKuGb0g/qO7n4ZFjH9cf18UnYG7qKZvchm65ow
T0qpY2YhdI4gntQRxoOS83Xf3FQjK6QzMxzAl0bc0vJMyrXEP9fGpjhrQwQQ4oDs
2TtvC51Dm8Zj4VOXpsGl09AkjNN7NIWTlvBw8mVoabL5tLBkShH+0GmdNsFr246n
ZSqpeoQb7fEj/oHBdO2x5Bmi/3xNeNZxhqbRmKL4yq63oPVKFtX3AVqSwXkgBegX
Eiqc/GP4COH+QluN+wY/HCDBVfi6Syz9PTKFC7Yv+xQ1lF0Y2t5X8QUKDHuuhy8A
WXKAEPholCzffGNyM9IX3ySNIZHx6xddxmJI36IOWwwP8k/BPkBOMIgULoJs1ecf
t+nl0bc6Ca6p5xhOh6M9FSFRiRhds7pouQWzQAbqwbmugiKTu4QgTHbGrLAE93sb
1f9Xerx7IViQhy1/XInj2mfV7Pns2uvVV01iJrJp6TRLI1qx6CKFzThua2Q96ha2
HTrQI8KEEBPua4Iz5xAJJd4IEhpAjisebuOkpleimAaxUT6WP/4gBjBOHFpIB35N
dTgYVB6bAAR2vjDKCTXNTK/TNwPmGV06DTiQP2vE5OvD+bz4Tss19eJHzpXdjJho
dudLekR2GPcysJtooMC0hdsyz0gWgRV4LAFO0T2Z9a2QxZCTS8ukF4YstLPb08ST
RWtfMXM936cY/Q+szud0clFLSlP6+8IU9pdy4GTPEQV1qYlv4ZVcbO62jFQl0ncx
eT9+xpJuiDvMUdKPnr27UL/ash/EpszUQhF8bQSKWpT03fgBm2rpHV5RvtXUY8+H
u96++UM077hkp+kcdbcMH4+xgzywPlR/vDjI5InHdGFY61VmqN5YojVomYuBbI1V
QIh02WfsUJceQOkMdghOw/kvNj3mISpWzCuAJ++st3I2F395X5tM1Mtx6cd8A6Sd
p+sZKC6puzJ/Nai92rUDNiLQq/aIPBaC6y6dFeOISDD3N3fg5WfF7H6Jw+dTe3FL
Qdubhef3oywOOZuZ9ecYzJ9Gu4sjNQVp3MnlT9hnI3a8YYkl0S0dwaIQTgBLJ11P
/jlNO6yiRGpjHm9vH143pvXxJLxXNZazQeUb/lUxa5b+6vhpTFWEqSDkVqtZyjsx
hKRwvGf7nkMat3tcXpnSlnVgQLRf6XyXP3P3iqOJzZUDENcQC8soMN33CnajNmdj
u3Rtaq+I+cmz+3fm1ow6URj+DZcPUR+7FmDR+6GS6OXZGKw8HNRRPvgp66olFq+U
EU1pq3OoUS4ZLKsjX7DuYIQyxpfyzCBAp9hnQ17agwWWz7H7fWEy/r/Bk3BrGvdt
XDN4P+Curq17XVlbx5t32qXA+kTvRRkgsYm1Bi9dZVBG24s8p4vl/sjzPIYzTAQN
1imiUeNOHKwLh9qZJ0G06ec7xSmei6s0zwLpLfDb889aTpzPlWJIqPRX2kWNrLx8
SHEHLcneNLdYCz15oo8I1nTh0waARxvBVO2uPmfF6LNmokVVe+1uljva1p0s5E7n
A2SeD43oTEpX5axIqZhVBStxN4jVpDrCeoHWAhXPwPj7ELjC5LSHuC54GOigERLm
m+qPHIDzzY7Ns983mFKxEznqbV1JqaJHaCBowXhtLYzQKCZSTD3Vpabp+eK3zSrE
T+YVDH3AdU53PBcdkU2/TuKWte03lPD2FC8GDw+NZ7SKrXK8WyMB04G3YXJMJvhB
2VKWHT2pPibBisTxZ6bb3O1+10xTb9wszqEaU4YBv44QXR08rFyPgp3eS1A6r28n
19mWzZMaS0J8iNzETHVuWgcXrSYuhft7cMdtnUeJfKfmnuVrAByFXae4zoLxpHZl
OLoV8cJRWLOVjqn54ecDVKT/emhx+6y/KX7GMZNu8kZIuQx/7utV0E9sHUZeWYVD
T3xK3pfB6rNyHD78jXjKaZoP16ewkqjRDZUQgdjW9hMkOd9RUrkW6sOvy5BgcYZk
0xzu2Xv81y0jEcXqX8S+SHpd87eSpeWWprRTFAby0SBaylqsjSBWwi6ClqIyZDq+
rWKckTI9n5ZB4xkDrO2+sECH3uiRdwhGFIKAuNZDn06ufHIZREKwnJDZZLCvkyGd
NiGmoYN4btiLSSE5uyU5l6XbsnWxzT17eDCySF592yiIfi0pqqqrpETtpKn3smIP
N4RzM60ZNU3QG6mpgKrpMSh91pplxwaRaKfazhbQMTJ604PoRHEwnXlJsnNUtQWW
gJ7iCYnqWf/Ecp+pRgm2X4CmifXxPwgqv71bum7iypg/Xm7HxllDV0S5S9vYzbKF
rIEOYaDm1ZeYKOorn1qCW64+9O1HrKQB0g4ag2tynowI+FTJJ0xSpHd92FBdrnhk
xPKM0o5BBA40GQkMjkKSET3+tRNT331hEhcFnULhwsSL8Z055E+T7ekgTR4xAV7M
Ry3UpSadwqk/yG8l1yxIWOT6oINcw/xFrLoqjkfwY9CUbAV6oDaBD5Ov11B6Mp5g
YfJgWUccOEtNM6ftLcTRM1GBqORhidsozBYRdE1feWSpVVDZctTUK4bsVp+/Pslp
oJa3sSt2bzJZZDehASpcZzSaT6NWzsmsFCCG+9Wc9OkQRL2lcKT08XS4DLmLi9XE
BSzbv2xSfobsQJIMCUJk3d4blSCOfk4ksxHnIwIiDmSO3Vm0MbTIu+JCL90nbj+6
WuhNZ/u9ZU+FnlV7uQeIyy0i3Fbyr68lHPcp7RrGvOh68hqfFm8HDY4HNq1lOLrH
J9sIHhxIMAIYY15XSe3GzCe0r0hBHytgLoROnSc5rBMmWe3y6P/uIYXFj9bTDghD
udwyHzq2lAP1rLYXsJZU7JXcKKU1D1OSxDVOJMBsK2BXl8iRdanpZyJKhwJS4otv
zwYAGnEMD6FUYKeUz9tz2H8ZvXBEgA1wYgqlXfJ5ilQEP/wtpitiRUsxvHk5IqNU
cMInpdiS3l/Dw1kYFIS+urn0ld998vQXrnzSqea3RUHpvbt9VChMpk6noOFGpHKO
LP6+tRX1zKHEpPoURQfLLbev+9CKfnKnUutArTHqp/luCC2nJdetwKoV7rBr2Oxi
8sbuqE8nz1FjT41EnbtyhUyMsIY679UupSUFFDKEbjxQUbLFkO3uDBPxgALATOLZ
CltlLCwy3lOxcBicqShYXN+YiBFu8fZrL52KK4irJXaFCDUlam2eP7et3Ezzy644
DIXWxdd1xdr4E/KCitEbkweuAFrigXbQgHUU0B+3QKU4bXrRvvCnD5ZTvyrpHZGg
Q6lLNp1L/LLxHRKl3sAmQcGDxNowWnqABraAtk5Vv5DTQprKz+FIX6n1rkvLJjmW
2lTNvtJVQyoU+/sKO1SIgAx2shXeu0/+XkQETtGV8YLe+2XG1PdAs8judT6ZvdPd
iXD2EcaKQkVtDq6Xp+6hXsJaFrw6IS4+1+iQyHjRuXxa9kENZkq3XtRVHWkG+mAx
IbTFEFCPJ9QVatB5OKVUkgTbclul9h6RpNKd3LnFZM2tXgnWK4QU4DupfLEFPFUP
4mV5/BmBBqjYuR26IFKHuFO80ybo1cBZmRWfjHJgoyVKf+dh3W0x0rU99kHy4Xgk
iVGgSF8fYA5gF48ZOGAlmcVDM7PM07t03XsiCwlXDFcWp+44Rztxf4/5Bmwsxi3z
3ulUOhJYKEdg2+f0IfGbFy2UNJdvbmqn7c4diw7rwfdTesmOot7utvj9sdO6J+Y3
Wsb6gG7Wxypb/7KpyKcf70LC0u1gbeCX0bkakHqlIk70n1W4gI4DkgargdI7BbEh
5QjRly+3Sr5llVzDmXQwzig9o+YOlOyiwWcuJA5Kf/1gEgFaCURrmb2rGXkeidLg
znwfcf/a3oGXC85cCy4U602Gp7LOcmwM44p9JQRFtGEfJ2YtCYYXYTn8C6elYfqz
NrjMHtlhDiwMrOJ7VGta93tRvTEK77MN+pzdvN0mOa8fSnVsDm4NN7u6hqviJ13C
Oy/jR/y7UMB+8Hq2Hvmr2SAMpmu4iswPwvfTLymnZjt92lT2ldGW5+v4Voe4iDwt
boBUHtr36Rqc2snZQvxq+Jub2CUAFZP/In4oHqodcbtqbyQFtnFRZiog4eYiEcw4
rjh+QixsPZSvr3VNFxZPXovyFtO2BK7j0XDjiddXqlNjjKf0CAOlt4hFiAIVxCLo
TRQk5enxh7ZqelMZCKHbMpcliwyCYYeBUcCXvoYDDpMZAUjlBRuKPvD4OBkWQIPD
gRjKziy1D3mokGz3hpZ5LBxFdEnLfKpVbRkwGlG1KbrqkqBkWmD1/YZaT9NK56V6
F2Up1RqDFP9z6kXybo7GG0IZ3Qn6X38RI68YVOVTXAWklXD8QF2lC/gCfufqPEiP
UcMy23nG69ywcKcape3kF8UWsFUze9VagV1nNhyIGtRtkyB3WV50E2YgwDofVhUu
o3VlWhKTFNqaNLQ3CILpyrHCe/N5HqRxddDg/TC2n25NKV0zQYfArpJuntpvgR2O
VA7RFEM5BphBHKo0ZsDM312Z9z5AyNyaumv2KIOPOPoBJDcNuiMks9IAHdGMZv0U
KXyacV3Fo6x5seoxbAQgYGTBtqbzgwWrahjSRQxGadXJkfz82q4rg6NQN36xVFy1
Rn5OlMk7Pri6H9gvwRmx3Gp9o5eT4xHUC2F6mrGrNddSGYrqGLW3fX/WLf7hJ8/K
wu2KBN0/moMpfmfBxxCAF7+MNRCSU2KyDIbYWS3Wh+SNORmJxWbUvm8xwon8Gfgx
9LKySxUvjHSOVq81puzReqYpq4hRyNEzm4KqqcotQRH4vDgrZOHYRyj9Zp7WeTqD
XNCctRj1TMnlEdQxleDvgeybWkA8FBXtKBpOpYdhcAKCHSMF0f6axbiUlrVAqhUk
QKwKfFYLi4TsT7JhXRZdsZGKghi9++kAla3HzcWYlUTlLgjSwVkAsZujHXYsFSx9
uS3pRyKG5FhufVRNhkQTxcr3an49sIs0af9yZIMJ0Y39DKkvgrjIA6x4GnRaxBjG
7W+8YhlpPfLnP8YcjkVjfZXpx9xtyQEXDT3c9rp6qTdkDoqR5rp2qAseDfQ2Tm9N
UTXFI1BahI8IYxgUH3PGF4egFOnXp/NSjXPA1XYpCIxX/4R/T6XgznA6YQIiT5PJ
Dg4yAOwEZc3FsIXWiL4bZL+Hpqs+3AhKWKahsFTlWu/FnMBY5Fo74IWSKHY8Docr
cEzAvKDFHCbKTI8/vk6ANpd313PNApMSmCsXG1vzojKIJZMI5sKwInxClp9oSW6Q
4GyF+3bajUXmFIH4aHEHLbwnfp7LpbWvVG6yb0v6oEr8U+lTcFzp/IWaouDq0eNJ
OVJy7O1PAdzlAdNSJKTe2PaVLhjqVBjM7y98e+ZiIDpAmvV/GvdLH7Z3J3Di6RZH
fojiTMZUv8IqikRakWssYfr8NSDXuP6AMuSfeFSpCYk+kBozOEOrEOJNuqmAnBjX
QCm0PMrq7MFO8m/k6B3IPCnlb9x6ZzXKUfZpROYF3pDSRuZ4xVaelYVEZ1EWWrdr
ITfkMldXfXlcURrKj4arc4VTZOev2yBCarz4zmU+9/O0AoexzWhvIicUGjqQ4ZLR
VMAjC8zRCH2tY+ahefBJBDMc6stT6OslGCvXDHG7tbv7GaIn9qfdKKdVjL9UozhU
F4aGdqPGmIAFMkFPMsjcD9ylB1e3WcCr4nzXUS8UoESmnIF11OsTROgW+RAhCH/y
Rj11sjEEwqlTp+ulZuwb+kQ/RUzyGD9xzL6la4kv+TlloG0dJSyAEKJi31+kBLvS
BVWv/FDdjppWLDcMFPUu2C8Ia7Didjus+JhId9QSRi5g4FgmOfGkTzkz/3oR4qeK
F6OQGuZIl76q79JES+38Y8WTn3bj4oCR7whL2tR9XFtFMvy+PmkZkfKhFDicCe5y
O+OMyx6biJCF71YKc+/rCc+JW5fr6uvXws973qPAM/ayaaqmo/0YkqGpc+Gp1s/i
G22CeBmnv3U4+0T28vNti8rMreqnfJhpKGJO5pbhAGwk6hUioyfLgrhlhZx4rMpE
YyqHZLDlMiTySLLnS9MCRjajcxS92qwVLbQat+RghskVn34iNoQ5EDYeyZDrh6Dd
Y7f/RFqYoM1ZkGW4rejx+5KwJthWVzjGIqNpino6vbfmVrDN34pePDAXwMe5Xtnl
VaGngvikuReE0pTfUQxV43rvgv8cAc9Y83LYdtDtQsrGasth3qTPYQT9A8Vpbbeu
rlD0YYj1trA9JM8X6cu0QF5qHWrH49mkwW8px0ftA3ovrZXckRfDh5geC5jtjTwK
MhDGsBEji5BiYjVqYUy8uN+QtrlOzWC4+MJqwf8/QvbcmJp3opGO9yfE9xaYgDuB
4jvMqp0EMxF+lXhKfZ7YcKFIX7NqkwyUIQzcG+84xip+7jDgdbqwaWpqxDrhblQU
ZkQSJiJMLvtuLHyxqwm+Z6geByCRdTCP33RPWcnyefxuSPlrfhSmkqH/mYmo3AOS
V6LHuoeFLUBoR9+/qCXxCt8IgaksWPzl3LMP9qwOIwXl5ZVsCOr/CIhKhm68P9bQ
ONl7q38L2wztEHc2ZZmJiTDE35lGmZhqRzpSwcAK2CPjoAl9C84neW3lWj0dsqYa
3ZNk4mXBF5tJY+GRiXplZHPvEdGf8lrc7vXccCVhz+wxvBVS4w/rWQrMOct0i8xe
OaModVSrM+LKtJqS/8Iu+8xfiG1uWxmu8QX/BAXap/MFaR5RhvQJLiGVqkrI8hJg
McVs7SvRaq4Mi2Yfh20p4vK/dRsbmhUquseNfGsLu59Elvh5UkUWAvhSO9I9Oo49
ng+LFQHf5tw8h/EIl9kOrxIk2+3iHiPiKwOPRrCnp6OvYr20Rycme7ZcxTT1aih7
/9xWtACLtEQkXABfR40TuMduIYUOLX3cSrhCYDvNIdOf/bvDDRicMROLy0uTdg5S
DR6zYHkyqwJIK7KYE8NuItw/YFK50fdgs8Tui07OpSw6BCuqsz7SzHZSyne6tJcA
x9qHTLdw+iSsohVldkWfKWXKXzJ1uS/47kOz8UVMAllabfH1J+DAmBG8WSJpG3Rd
9jq9gTZa2w/hnK/FhrrJpIxpS9RW/cj7sft8vYMu9QoagIIFas1olNjcWTViDJ2q
sTgvtb/HZn8elL9Gp6dJK9Nb1WDAn6BuHkXkNV8FGWV/1amTMl4nItjuEadnojhb
b7P0urVbYzMvvxbCiTtj6Br48VITMfWQt5saNr039HzHUazFSZRx3aDsirIsv+m7
CDDVLZO4qlizmB/TveTp291BgVF7ub/lHYZmR5zS82jysewN8okf8IQVzLflXQik
RzCSf+LWRIMgaC/lCcheoui5PnIyHZdgiQD2+jehovi9IuvbwmwOoKuemRvw3cun
saXCdESpNVL9MjSr7fDG4S7wdKGKnnBfNmx7yxAG92SjOmhvG+96yf/S2rNluD6K
VDebemDCD6qwoN/hbDHPhLgCkIPn6JA9Q9XJJRrHLncilWTNKPoJuaNhDjx8eT5Q
BZHqK7efuRTNcPbgtsFuTVKphFvZIFlvZ0/bTh0brxOOBXLJaOZRZ5m4Ko/68GlC
/IY3eymAu0jrE2PFWGEDq5YZbxB7xpuWz3cMoVlo/SIayj/QNEFAMgSiCac3IUYt
MHawVh2K+Q3Yz4EFWfUHhvckv9wB39bIIBsgtnvqhozTZQMcLr5F1UHVHbp6g5OA
TJvUOfZ+9lgFMQNdsje/8Wa2eQ7FWpXVudtYeFWPPeaGHGc13q/htS4hp5GD84z2
tsMTbau6oQqeQKIxZfvzBESmBX8UY2fylMvHB2+cH/RjIOkKuGilnthjBTUqKnMU
lmdlobd4qarFwPkECV5Z6rmSSSMsmCRsu+XKyLKDO8Pwgq6Qfm0xs0tRIpacjGTL
ezxOfueiiVd0HEFsyp0dFWXb/hDwTcZ+ZqEYnqkKWjieq0inaSCBD13E7QAV+brF
Yq9r5o+FAzS2HXNCJavk6rVbfLDoqVqW1nyFWMy4263O0gNJES6pGD/nNhngwxIb
pR9vkjo8t0f/j5lJ128wJ1LJqQGApB7skDcU4IqW7L0WDPLwujRpySjFIxd64Fsa
2nUY7vOYlp+4LIdqBmfx9oLXvyHAcu1YdyGjpbgzhVzLOcIN2TFUAcBbd7hrFPV1
3OmnD/t9OLiVEhLiOGKhUj3FGugMFFjTtJ1XvgurDTY1G6PSlcM/I7gbhqOqPQHp
2WvhhchSiOR5eQpI0VwAOaZ1FVCzuj4MQX5m6QjxvheOxj4DcawzC2eU5NPpMfD9
3SGeN6E5O6uf1kIGIPW2CPYn36sijq/uo3J9/pVY7UJjSmHZR9HggTul/1usv+pO
cvDNseQRgZrKvy/UIocpcv2T4oyAQbeYp1DJbY7I3mmST/j9E3w+7u22upbWeDcg
N5efejqAg+w1id/jinDvFb4Tve8k2VatLcvnbCY8hgAgHDkTCrBdherQ3sKGT4/A
k61xxWWGf+YYvVfE8yb9FziaonKaVqw4oBvJ5Q9KKDF5cW/r+oCMD6/RBSsANCHC
JMbrqOGM0IeOhPEAxJUcswdKoMQLh3rVcQ4mLbGyc+qT0Y2nnqQ5Egu7dtWdYMCu
AlsG1kzOaKVJYydXbG0jFy9vmL/lteTIU05D34peudHB/rV/cbB7PFOgVNruUcEC
dPhAaKscUtqo7bP8sJ0BwxTTeyrRy25isBA55iJAUXEGa6v0xtMSO+tFhbGcAucM
mBxXkTuJxCq6I0Q8x/4C9y2bxHWDPCHAA8N7wVSkGPIn0+cPxKgfeucnpNnMIerA
kOkHD4f3lWxlaNOFpQ601XUiBH2QcjS6H8/c9ORXPRc9DwxCy+NXWGjpilYj+jRV
Ilf4d99yyTKkpi9ADazfbeB5tWhm+RpW594SSPS025q42b/q6NuGo4gIH1GT+tsI
dO8Zo1vi2ykRiiPgGl/CNFRYyaC4pUN/gGw/LmX9mbgu0A2dicuzsW1OYz2zFFSJ
Ox/Js7EUKAxQtNWMsp8Vf5Xrkw/ZSLkRVRE83qvcw1u7rJGpdzi8pkYehvdtKQdN
CReCOUijkI9l97KCy6pqp745JxKjlTHB6IzxTl3EnOGYo5jLLCsUf7tmaXuQVfsJ
fnVe+8XK1KS2ZI6lTEhvPlBEngWPfHrpe9Oj8TnBKVSMQeFQAC1j4V1c+wtkCCrq
DfK77CR6soCJSyxnBDfsFmRJ+w3ze+bm2eWk3ZbjB8MC8nsSjbmHo2/C9fHw1MUP
oNj2Y8h82A9GM6rmMPm5Y2hqXV3KpHk9vw/7z1S2rNUc/I17kEfnmT/hBFdcazl1
ksC/qIlykvhG5BaQEPMHjKra8c4ILEVgb/U6xNNf4wITwhqMyHD9ZvoGUlmiPNnQ
e/ZHByfWgQiK7Gops325Dyci0JQeeX35Gfi8oAVVC023iLltfYCFqtcIgAe6uhNe
/5CzHo6k/+tH5D8HObzoAVREIZuIbdktQ2KtsmSAotyQHZfwh9y3hxlnjqMkgjak
90rbyCxv+XRVL3lJzkvxMlBhJPg1aRc0t+q8GI4JzbVeZCtOYDAlnkdVa1AzB3cr
JXibWG7Qa+SYeLTJ/4B8HZxyH1jIdnm7L4nOMw2tHI5uJ6A0LAnxsYNrLfZ4MtRY
TlbJTOTRNRqqSgtI1iV9Xzc0WSSB/JnThOumNeUceA5obxPzOOedIGRzJ7h7oVyN
1rOgniOUvLMAn4Hvx/gQ/D42Cc8KB9chY/6/BMMW/d6IbTsitR3+pLWiA1EIKa3W
CUdNe/GKBmkMtBQVZAkUvxg9bm7dlXjp4wijqiUcuGOWF2qgj28eIe1TiJIq4OXr
dd/zTxK904r0bCUZJmWa6UCgMMzBc8PyWRpssjXlKygBMvrwTNjwYswjlS1X5R6S
+9yQ2F9+bLhjIt/0sZmov9GeYJySedl2vxdSuovLJz9RmPnLcXHiwnB75pnmv0Qx
e8WJ8AVaaTXcnndrBMj1beymdcAbHlzXlVKFXD2uU25dM+Vgwm4HpZDT34W5AqXj
7bdXLv0eU/PO135p37VosVBwKLFSj/PAXJ6BM0bcgMwIuL9qSKvoe13CcqruMVCi
OwZMl7qOHy+vxuX/gzhcWt34YC0JDpQhKGxW7Iy1sOOKbFjFoZsqaQWcqX5wGL9f
cj+bsqrKQJfWikN5lUMv18kILRfwXG6opWmC6Z/3gnnXC8AWEnqicLNhYXPDZRTd
f+xXomld9Jl9DCMwJZfofud7IkQoMiJumbSrhTY6wH7APHYcIIcekC8JEsVE5BYd
VXkBu60YFFvhGDcDNHdfZnMgGMMTh5VAi+p7duUdYAwMd+Wvtbf7+CFCh+x66Aea
cuOmQb/OJnz73jito1rbolSdypWJoNJpzEza/llKpGkxxsHSk9wD2Skm+MiIeDjt
R4owKOrkFrhJ0mIqGP9bzaVqEQT8wFnaElr3EuqKS9R/jN3xVol0ZgQCFA0GyzMX
Gk6sO7F7aLNyLwug8NiGKpjw8OEB+vb359ADyosK4zIjViGT/9K5xY+GKUyNq8Oq
0vj8AkjYcofaXRXRjj8iNGA8QmW52MxCmn5GeBenyCDoPUvhGpOFSSop3Yn2fFo5
DJNcX5tGCQri45AYvIDmiLpA7gAWI/QWWzd45acQJZn2f+op0PdcW+SB9AcqMZXv
LdpocR5ZT20YPtVXnYStHDS7OzFGDOWVQeoUkdvu+Y4aYOm4Kn0ybx6PxS7llhOf
GQckcF/l9JAXNl0iFdjkSRNjpTMr5oMXD2ILr4CzE9GVgJUV3lmgKhFW+JV/EtY4
SIj0wlImhx1sY3WbEm9G/OdKqZf6H1p9dEENtFB8V2QQIoJXNQcR1RzmkAyq3XOj
r/f2Ak5gTq0R3ORYeQnhgeEsNLEZz5CJZMJf65e1U5ROzE191j0K+PHxOy+zA525
iwAXYO0GGDDVXd4tdxPsnxw8YDEaQxYaJNUc8TUX7faPQ39SU67ZzHO9caKpHVcu
q0jVfEQjL9rKO0eK7eLORtq8dvxRlQfZ9AubbN8sf3rKeZQRLO8bEj51Jui+b6Pm
+9RJCDcAdf7e5GMubvhIkAsvrbBObp0Ly/dfqbh1woWTYXn3hZo6ftCMepqcDw44
b6HYWmYyWXHHvxsv7yuQe21ihqorevxj3Ffxe2GcNnxjzz2JNvuK0h3+QM0dnfts
BvdRU04OhvE0M2FI1ipcvJG5NGw1dv/MxUeCExFadrxfz8HiWAfP8RpBeN+nOzj2
PiD1pZms48C3PtheEGLlfSfJdMBTp73j4Wl7NNNNBkME+RoUgbCFKdDeCpcwPVCZ
f/blUZl1IDJqkfsrSt7xaA==
`pragma protect end_protected
