sync_sync_in_altiobuf_inst : sync_sync_in_altiobuf PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig
	);
