LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.ALL;

ENTITY DOUBLE_DABBLE_8BIT IS
	PORT (
		CLK : IN STD_LOGIC;
		RST : IN STD_LOGIC;
		DD_ENABLE : IN STD_LOGIC;
		DD_IDLE : OUT STD_LOGIC;
		DD_CLEAR : IN STD_LOGIC;
		DD_INTEGER_IN : IN UNSIGNED(7 DOWNTO 0);
		DD_BCD2_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		DD_BCD1_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		DD_BCD0_OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ENTITY DOUBLE_DABBLE_8BIT;

ARCHITECTURE BEHAVIOUR OF DOUBLE_DABBLE_8BIT IS

	CONSTANT DD_SUM : UNSIGNED(3 DOWNTO 0) := "0011";
	CONSTANT DD_COMPARE : UNSIGNED(3 DOWNTO 0) := "0101";
	
	TYPE DD_STATE_MACHINE IS (
		S_STANDBY,
		S_WORKING
	);
	SIGNAL STATE_MACHINE : DD_STATE_MACHINE := S_STANDBY;
	
	BEGIN
	
		GLOBAL : PROCESS (CLK, RST) IS
			VARIABLE DD_COUNTER : UNSIGNED(3 DOWNTO 0) := (OTHERS => '0');
			VARIABLE DD_WORK : UNSIGNED(19 DOWNTO 0) := (OTHERS => '1');
		BEGIN
			IF (RST = '1') THEN
				DD_WORK := (OTHERS => '0');
				DD_IDLE <= '1';
				DD_BCD2_OUT <= (OTHERS => '0');
				DD_BCD1_OUT <= (OTHERS => '0');
				DD_BCD0_OUT <= (OTHERS => '0');
				DD_COUNTER := X"0";
				STATE_MACHINE <= S_STANDBY;
			ELSIF (RISING_EDGE(CLK)) THEN
				IF (DD_CLEAR = '1') THEN
					DD_WORK := (OTHERS => '0');
					DD_IDLE <= '1';
					DD_BCD2_OUT <= (OTHERS => '0');
					DD_BCD1_OUT <= (OTHERS => '0');
					DD_BCD0_OUT <= (OTHERS => '0');
					DD_COUNTER := X"0";
					STATE_MACHINE <= S_STANDBY;
				ELSE
					CASE STATE_MACHINE IS
					
						WHEN S_STANDBY =>
							DD_WORK := (OTHERS => '0');
							DD_IDLE <= '1';
							IF (DD_ENABLE = '1') THEN
								DD_IDLE <= '0';
								DD_COUNTER := X"0";
								DD_WORK(19 DOWNTO 8) := (OTHERS => '0');
								DD_WORK(7 DOWNTO 0) := DD_INTEGER_IN;
								STATE_MACHINE <= S_WORKING;
							ELSE
								STATE_MACHINE <= S_STANDBY;
							END IF;
						
						WHEN S_WORKING =>
							IF (DD_COUNTER < 7) THEN
								DD_WORK := SHIFT_LEFT(DD_WORK,1);
								IF (DD_WORK(19 DOWNTO 16) >= DD_COMPARE) THEN
									DD_WORK(19 DOWNTO 16) := DD_WORK(19 DOWNTO 16) + DD_SUM;
								END IF;
								IF (DD_WORK(15 DOWNTO 12) >= DD_COMPARE) THEN
									DD_WORK(15 DOWNTO 12) := DD_WORK(15 DOWNTO 12) + DD_SUM;
								END IF;
								IF (DD_WORK(11 DOWNTO 8) >= DD_COMPARE) THEN
									DD_WORK(11 DOWNTO 8) := DD_WORK(11 DOWNTO 8) + DD_SUM;
								END IF;
								DD_COUNTER := DD_COUNTER + 1;
								STATE_MACHINE <= S_WORKING;
							
							ELSIF (DD_COUNTER = 7) THEN
								DD_WORK := SHIFT_LEFT(DD_WORK,1);
								DD_COUNTER := DD_COUNTER + 1;
								STATE_MACHINE <= S_WORKING;
							ELSE
								DD_IDLE <= '1';
								DD_BCD2_OUT <= STD_LOGIC_VECTOR(DD_WORK(19 DOWNTO 16));
								DD_BCD1_OUT <= STD_LOGIC_VECTOR(DD_WORK(15 DOWNTO 12));
								DD_BCD0_OUT <= STD_LOGIC_VECTOR(DD_WORK(11 DOWNTO 8));
								STATE_MACHINE <= S_STANDBY;
							END IF;
					END CASE;
				END IF;
			END IF;
		END PROCESS GLOBAL;
	
END BEHAVIOUR;