package rmap_initiator_pkg is
	
end package rmap_initiator_pkg;

package body rmap_initiator_pkg is
	
end package body rmap_initiator_pkg;
