spwc_spw_tx_altlvds_tx_inst : spwc_spw_tx_altlvds_tx PORT MAP (
		tx_in	 => tx_in_sig,
		tx_out	 => tx_out_sig
	);
