package rmap_target_register_pkg is
	
end package rmap_target_register_pkg;

package body rmap_target_register_pkg is
	
end package body rmap_target_register_pkg;
