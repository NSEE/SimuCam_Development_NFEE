library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rmap_target_codec_write_ent is
	port(
		clk : in std_logic;
		rst : in std_logic
	);
end entity rmap_target_codec_write_ent;

architecture RTL of rmap_target_codec_write_ent is
	
begin

end architecture RTL;
