// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
FQu9f41q/bFdV6gRIGTus5uv9z0z0ysxiM9UcAhf/vnYFcC8nJQlOw4J3b3ubEDX9hJFDa6Fa9jD
bZ3emKazT8/DtRzlNHpAK/32nDzGhvjefyxK3njBRsA186aSYE/iaGAcVizvb7o9DvlHemG02Zo6
XhYbLOiMrTW+0YKvf4uecLGW+Lw+L4DGqt2U36FB8PXHaoEENxTD/zclFg7tldPoFPXL6rqMlZfn
KDEclrifwytM0qHEziehN5Eb7rim998EXKrPzbeN4Is23/BL3WIUJrGFtKPXyEvoDG4YAM75TeTo
E2IB2sdt9qVekHaLKMZtgHQTdLRNeHvrhHpbVw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5264)
nw2Bw5QkzY6+AuPwz2hGaCLvYTQtN3U9AhbVLX3de9fePn4iGb4NJPeXUR8/5+nBZMeaE9tUWroh
9oNqcyRZ5iBdQedX6ZDZ3tLP2Kc50a55oj+NQ2n12d0ZnVABl9ylFu3mhBmBQAqXvvBRZ8lZ3PHM
9WS/1tjD3jAfL0nI6mbUCvSD3B2tpnI/mBdWEZF4pUYy65jaPFL6GNpVrFk1VBA3ZcZLDji01TYt
IITW2GI4APCvSxuXI8JPh85+VkJW2s0rb530YI4l+U2Yt5TistjCFPUcaDyiOWpmNiexFKyl8ttO
yfIyOPoLfAGz9D/8TbMK2tOc0mGIl8XIBp4/24FKWNVK4JJ4fbJaL5+dU9IwF/5xZKqRKIM1S4dT
NMI9oeIRmIuUnceNM9pbL4lUQyngK2unbfyoWgLEo/sk1D7cUEa7GGmQW1BX3Yd64pGv/cAx2Zxn
s7K2uejLCHNmZTFveKzq4VkzOAjhdZKSygWtTccX5Ina+xVApfIN2XETQY8wlo7IONk53KsP/S3G
z/BktMBWxfgahSCync0nMYEZI2Rmy1NHK4or0uqrpWDiWEpQixV0N+NtC08fMJIScINuIyY+7mY0
JaO6MHfziklI6+DxLwvhAUM7/w7NqBusr4/Gzt+kCDaaQThINuYXW7WOZRuUpo4kkgi28YCovM+q
ts3d2YxFTjW3RuyfGRNM66eAMcvFBZItV/NR0HSybE8CTB9V6tEISXiAw+UGrOCEvcga4w24yQO0
8XZKXyvUc3bTUSv3+/JfUtorOe/pkSwoGRM77aMUvLVu9cl5Kj0QsHyRxI6qvLJc8fxp+SH3z60e
lklQVlje2pSq5KGpnLSvOBy4rVzDQPAVPyqLXDby7qVZ/LxEttaiOUISoVIuCatNIjzUt+L2fnm7
uoXZ8L2U/zAhy1kQJp+HrFph0K+p3AWAxP5oKAQolMxk7tSx7mKslB/k6EjsRaC62aTBIIsCeh2F
Ftbcv+0FiH60xMEYeo78rksnB1sSEP0CAg+ssTh0vMbJbi896+u74PSwbKEcNwp4hoKCex1TzQP4
XackYlMxOHe74l4CYY9f3r/oPaUiHZoKe0qoBLmIqGb0RGvg0MNepblztGzClF0LHRweDa1XppqQ
exnrYpe02v49oQERFX3+CZ036wfzFRWzbHXsEx31Zdwq7KGmaAxt+8JFOwZFc403H+QNP9zCi37Z
jd8Gf/Rei3xGuzpEWvqqul8LrY4kp5HZmDH0Du/T2A+H91eoeW5N+TtJhxLE4M4SKeVIpTTopQI/
RE9y87rjb1oo3inMQFNYlC92COwNhy4nr1FgdZ1bQn9x6IE6fYFRaubPmkMqw3YZlaZsiIgzR/Ld
tRX4XQyp4MxPyx92W6ZULqXKIF6u6BssdV+g+ncC+iq/2LWRvhCBzFdJ7ZD1RBm5Q6U0Noa04Y/Q
0r3RE8PqJSbfbx7V3piNunc8VVoXUSDzcdHiyVIbSoIdmkeW+m0zF6KiVwoTsMM2VNc+YEJDuSOU
0wtJsVvL78o4pE34x0prLM//FqHAeIZ7bYQrgNt2VYAleb17rDkrOINP7HsqRmQnR97/peD+epKJ
kBrp1v5Gh/oQ0ngFxvOfC1/jRVZ7JTPjX5fbN/lUHJuPuMkprsx82egsRL1ipcIuWmpryPAiUyUD
Ul37Gb+nIuHJ1im0YOU5lZ66szFkLZakLsvPmco/VFRxgZxs/5SqLMRygA8hEFp5xsoamv7WbJ0D
MHNsO6KdpF4+yOkOta4Q1S/i1T7yFJUS8SuyjV5L16nYqYnqnXjTHTF95ctskqPhZHBy7yco8PRT
u7lEyOi3DwwC5Nd9ju/B1oVxDSQu4HA1JYcvl2+K6a0mxmSPcYPykrYHhrpJHiR5pudm/W87QofY
OsB9CS9+o8ost6PpBYMUbX4q53fsrmD0sL7E2spwdUTCACvh1GprgBrpkDm3DrE7LJSqaQ4sVo1W
1v14uVDqdkAEJmG2TFhoRvWp4Pb/7UJ5omLGlQGnwrieRuveao4sc7BbG7V2Gl7WUU7OugzAM+gJ
eBFw5jHE/NGnPL4rKaCJbSgo1Si31ezIBYfV/He0WEcFsC1P5Gxuw/pxCgNCHBhxKYw5sF6F235W
wFXvecNX7Ap0brLb7bl/HGDCBElj30EOdpH3jacdxFsTj1+0Aw7OKw2Rtt77BURfam8EuNK+db/H
4uJ58jSyptjXXjbyNt7c3aLEeX20IGcqYZqTNdd+O0IUC6HsgBHo/FMIkgOHhZJK2Xk6ZdCYUnsL
XgtT/e1lnlAfr8rnZUY2qtl3qxHJNMKgbueSjgDtBz1nxpRVY+s/pYqhFIGFkpQ7L8YBrXbpjywL
fmd5LzNewb49ki+vrgLCsd2TUxj9ekAD6CetmZ8WyBdzQdI+6ukXOv44IHEDU+DGV2KFvUrEEqEK
f9geCuoivEKtx8QFKW7tBwbSvCHfRlgL0s7A0mQ1gGDzHE88xUlt050roZ+vnjzFgwBBGIYVAmex
2I/YR9BmqjY3jgPt622LtcI6HXN6RcT9X12SZVlxmUqhNm79mZxZKruNBtIjFcprLCDJUpy7novU
4ovL5M9xyOryvuy7wR3gS8uvEegwbinT2t0Sb9vcetDMsG0siWKwXZmTEZGvpBmq/sf7tnxahkdH
8WZOyTVHNAdOjGHExVtsvR3O3xAX1XN6iGWndtAN4ja+9tkT6nEdFYM8flteLsbIKGKV7oUBn/a8
zBtrXBM6l+iWBxmCKJIyMyjVVFVSO6Gk7fRSV5TOWc9VdmxshUVZDToHG1v5Q340Ymw8qYXOaRgG
/c/xvWgH9/HCsMnBFKAmAfxMD+BEZcpwki73sBA5VrDnBzGM86MsLsAKhEmmah18YDx5o3127NU7
0ITZp3iIp8gVztnLJ40KLHJRXsfox57imOq0G36sieiUFFOV2WjqpRBIalTJoElXfMkkviqQ76a2
THButO/Qmb+MOcyCG/hHgOuTAyXYzoIx3bgB+ABlPfTwsp0OeaJJqBrUuvYqAD5RT6TGm9tP0XGX
NikNMTPutSKg477f15n39AuFhqAc7JGgXTM0udjMI2nc7uzIvuYZ6iK+I9YHkMT+lzzQ9vnDBTUu
WxtmMwB6rpYmE0SB28wsEzRYWxHPVegbSE2K6fimkTuYlmmeHuiSx9664fHdNHkSbNvrkbLt1REe
GsXcG7vLjNMfI4z8NcD9Gn46NYJ0NcuyOFAsXOyzdVR8tIPmDrp/wSaTcQArE26IM9K4dvLUyEFg
k0T6cFjTQ/XU5pYVBfdddejhePY5GbGhHK3QyEXY8OnXqgFATXnAdx/JX4nVop8etYzDLMaMxMSz
W+wmfQKcjmhV+7frBOEGSO1VrzGrbMskNRCgBh8yaTGk8Vz8xGYZYbnocPuEYZMP7CB7ghy65M83
Us/cER1P+RgMu6Z/NCb4tOG/pes2VHWCpixGX0wPZNrNv4Z/vB0RMbBApAhtFpHjPDd3H/rhiu49
M2aEewAx6Pib0gj7lgetV+WQB+NdYQVh+ZlXhN9tQldueX5nH29X7jZDSaHGpU/1X5nY/eSYPMVS
vj4nTpsu50O0LYVTqVeAp1rh0hIeqFM++zaRbGw7DaF0uyMuUidA36+XYaBog9XGnTVlhONhaIeU
/Q60M8yXlnv2vbqRWA5W/Wo19OLvPWmfvWcriR8Xy0/41tVagoFMhkUjbnP+NdNAg05YGfqrZHjy
H5EBdbouVhU7o3T7poTjHPAcM/T9ZWUmaCFkcd5JT8CEkhAN3YueyEOu1qSxB6//vkVCpxI/25ME
6OeR2qXkDtsOQNs1GGqmkD8IVD+CnubHkuzm94seHtn79ENLlqYGgoo6eV1oDpO8209INwLKQqmJ
SrgNa5IEb3uzycRXJfk92w0JX9ZGICZ9X+grDJBIjW+v+lC/vqB0Y+TA/UTR1fPWQfSuV8rY6VS1
oo2aiaIwOatXouVpRNfKx7T0T9p1yO+H29tUqjaTwnUD2SXBnA2ccmsJk0ceTFIBLdMPp2tgFdJP
V22XOrRVFlpoWAQo0TaVTu2bS3M39DJ/xfPRMLuKer6Ihik4QduhO+kP5G59ey056+U1s8g0rBka
7yyPfBj9GE9PT7z7zjQJi+7YDTNu6ZI3PGP23C7eeumQDxERG0ywaX/olngK5gW1Vl9/tF06NW22
KdJOr1N1+kN5X3seEa7Lad3hAoxL6h3SjR9wS3q4or47NCRy8hNHN/75BSl9XX4+WA8r/jEWpQkH
LpoNHdREsNToElPXB/iDWgaeoxO9MyaY0O10Mow98tfBz06UA6kHnGy7Nx08VrGtQl6P7xNjx9lZ
XZ20+zWR8KrD4NMRaUVjl/bFK+EcKuCxAEGN/K/8WVVZnEzdaQ47Z4izs8CCVWbny4VQK1a766FC
aEgdifJ1iI3FhaHHF/OzXWr9+nOLEovI7EGTyltRvdryQI/fkbZ8XLmlmjZsa12C8lI9Aa5rT/OQ
dR8e5wvj5y3esms3lFvPj0lLcpjVEY6d4IDsbkEAgCZnEnUquadxkrBmwD2z2H27RhBFcTvjL1Gr
Z01lHbiCS3hDCHWZc87ho9Ubn+q3dE8+OzwT/nhtkb8B8T/QpF6Xs3R9eCFtPMWQn2H6LbWcqsBK
UD5sKtxKT/EsLCAieCj6p3tWd9CRgevjrNcPgBAzbbMe8IXkOls2D/YcxvTmebTKulPDLPozGkb/
fy+5dzhNhcrn88xkb6zvBORYuj8k/Zm1+q7avVV2WyfuRtfN71mouxMb7Dicgs8YRYAF1sqMoMkr
B7eQaNHYqNmfCuQVUgb1UHxEIIGhvsirqYj/sYg1SPnMscRTE8jIYzFGojWHdlC5CccPupaVt61G
vye75IfLI9vAY9s8lgqFX7njvUgIirS/Jis8L4OGszK05AVA7iTfho/aASPU+ICwLV8JqKZ5dEgU
eYVEwc2bbRU/haqN+mor+VhLZEFUJ31yfnubtcuLmRZHIDiGMz+h1OuU8MddSFwuiXEtTcPUqfCe
fas5siP573xqIdy7pduvrsbgvwiaVnHxD9vynyZlrEHyorOGSlEav2N1IvmZ2Ix3d5usMP/ih0L6
dLQI8gTtOckOuG5EcJFHvMoEpHL4AeyoHhVz7Yt+nMDD5zWOTBarMSYSB17g75rFNpv9tBdS8MSf
aG6yD8lLd3qi2rkzM9Qoc1enAZEXm5ZQlA2P1M0BYIiOFCdDimOjgPOkEEbXIeHL1KU6kDDKrLX9
rzOgSvIYbi5lzROaZOit31GmxYcril/YkVfR8Wvhg9x8GP0KH/z7kEmi6LSK2ePsDM4vdRmyCxta
53eYss1YU+FJdcmGcEVjGThhc91vPjZn+DgL8kmarOrOhpbZ5TiQr+Gb5R47QFPegkyy6Fct9OnR
+lZmWEfRXF8y7aoP4aQOpXH99AofsejvhZuMw6nl5OQVKVc9Gfp/AxwRXEmXFjFRKSdGmRitw/0U
EkPGUAuMyqW8DkjrRhG9Go35CCAqqdMrEc60LvPxBGfic1EMC0A1izlpST71ulBBrV10MR3oTtZZ
EeCrz0CL/EkKT6KuA3aISDBe5CmDIyh9YphCt07IZEa+a5RPWxhcMpVR+buf4dxsRxf55woBfAEc
bUfu77MHMzuSorUKjBBRwNZql9l6Dl8q/PQnoY4ZymltAD5R4K6Ow1vl2mkgiIVxEYz7Y3R0kgs/
INav/O9GSssUcgBXzlmU8RIPhdltqobRuE9laQi/ovKBOw4cdZgdE/2Hp1DoKIP+ass9iTJEUStz
L1YnGwyYt0REX5y7svVCOXlZVuo562HImgSdxm0+b2xvgBhmrUReRs1A4nNJ+Txi5r1bGzsrxsDO
t4j5zsw7+w+ticEK3xTMPu2+Cgv84CW5Bsalc8C7gVbJxrDm2waOi8fF9RXh+KXRpzmXM3MDZIIk
kZrmBWS2zI3tIAP0YWheXkshPSZ3Q5PIo0RjCor6LHg5qW19hV3bKRxTd2Wp18gx4TcCNbamBAaV
HPWBvxnljDvir/RHBb8CNz3JuIZGInGaF7AfjIOnVgTqRB90iZuv/tjkdhfBe11aX25omnIv2AzN
cie0PuzbvovwHH6hMPKSMWYsQ7IlWrYkgBsJWTwxmbPDkmU5UiicOqzohRQSQfor+Wtnhhvns4gT
7v7xfxc4AdcTp4sT73zgmz60gFkYYTV6MUdmQeOS0ftK1G0Smv4Hb8sxD4hdDvUwwknuyWfY6zGX
TQp5ccx2UtMOJhdPREaHaOAXOI31alTQ74FZMbpplEjGTy4e2TKQh1yLeSSKiZo0RsTikLsNVpgj
QEx/k1vrOcbpyunuP4SuQsu/06XufWukSMBEI5+qTy9oUrlpbtBgAmGbJ3+ZCBYNIt5Z1lQXaf0N
T6Ume7c2DS/WejSvS6t+KLLZ3Es6VtbXMSHznI9U4UW57ju0BNZ56mtfFPo05wfS7xM354URDs9W
WAYPyQUMUDs2nWPNa+FM5nQO+o//l/TTPoBASKbY6QijZLmX7aTFRXEjSSCwh134yBo/dmKdaywJ
22zpXkEyY9goc9KezStbLTgAZzO+hdfM/3OASOIpBB0E8U6fZKes0cz0zj1NbnjwucvLJCvKa0DC
/2zlwPefS39m4HtGE8cP3/hM1Moz6JRFP3PsZW5DXRjOwBK3pe+tg1ZU2pMuOLOulsbJft2k7H+n
rDWawOwin5ndkrQgmGxcR8NTE3XnS7iuDY9BejX3QIWT1Nd5azgj1hC3LZduNZw4AT3Apuz2YTTt
zuY0gaIYCZFuxD5ufNqdVs90xDRuzRtj/GLLfpsPdFEw6DijTQgUae/VvM/st8OLGFwo+utJXHUq
tO/i4WfAIqRqyEFz6LAKsUymRehiRtjfOl1lk940m1Y8149+89zOmAV5CRlBB17Euz0BI8QbB/G2
ValVAMT3yumfxYbFqzUKNPP4da0bHwU2qUbzOA1IwzdzGVJfVyUX0C8PpcCYUnsYIa/mN3zoAbm5
UcLUSsYfqbWzey/XXB3RQZOVas0=
`pragma protect end_protected
