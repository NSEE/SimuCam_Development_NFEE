-- dummy file (placeholder)