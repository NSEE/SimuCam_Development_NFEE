-- MebX_Qsys_Project_tb.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity MebX_Qsys_Project_tb is
end entity MebX_Qsys_Project_tb;

architecture rtl of MebX_Qsys_Project_tb is
	component MebX_Qsys_Project is
		port (
			button_export                                        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			clk50_clk                                            : in    std_logic                     := 'X';             -- clk
			csense_adc_fo_export                                 : out   std_logic;                                        -- export
			csense_cs_n_export                                   : out   std_logic_vector(1 downto 0);                     -- export
			csense_sck_export                                    : out   std_logic;                                        -- export
			csense_sdi_export                                    : out   std_logic;                                        -- export
			csense_sdo_export                                    : in    std_logic                     := 'X';             -- export
			dip_export                                           : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			eth_rst_export                                       : out   std_logic;                                        -- export
			ext_export                                           : in    std_logic                     := 'X';             -- export
			led_de4_export                                       : out   std_logic_vector(7 downto 0);                     -- export
			led_painel_export                                    : out   std_logic_vector(12 downto 0);                    -- export
			m1_ddr2_i2c_scl_export                               : out   std_logic;                                        -- export
			m1_ddr2_i2c_sda_export                               : inout std_logic                     := 'X';             -- export
			m1_ddr2_memory_mem_a                                 : out   std_logic_vector(13 downto 0);                    -- mem_a
			m1_ddr2_memory_mem_ba                                : out   std_logic_vector(2 downto 0);                     -- mem_ba
			m1_ddr2_memory_mem_ck                                : out   std_logic_vector(1 downto 0);                     -- mem_ck
			m1_ddr2_memory_mem_ck_n                              : out   std_logic_vector(1 downto 0);                     -- mem_ck_n
			m1_ddr2_memory_mem_cke                               : out   std_logic_vector(0 downto 0);                     -- mem_cke
			m1_ddr2_memory_mem_cs_n                              : out   std_logic_vector(0 downto 0);                     -- mem_cs_n
			m1_ddr2_memory_mem_dm                                : out   std_logic_vector(7 downto 0);                     -- mem_dm
			m1_ddr2_memory_mem_ras_n                             : out   std_logic_vector(0 downto 0);                     -- mem_ras_n
			m1_ddr2_memory_mem_cas_n                             : out   std_logic_vector(0 downto 0);                     -- mem_cas_n
			m1_ddr2_memory_mem_we_n                              : out   std_logic_vector(0 downto 0);                     -- mem_we_n
			m1_ddr2_memory_mem_dq                                : inout std_logic_vector(63 downto 0) := (others => 'X'); -- mem_dq
			m1_ddr2_memory_mem_dqs                               : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dqs
			m1_ddr2_memory_mem_dqs_n                             : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dqs_n
			m1_ddr2_memory_mem_odt                               : out   std_logic_vector(0 downto 0);                     -- mem_odt
			m1_ddr2_memory_pll_ref_clk_clk                       : in    std_logic                     := 'X';             -- clk
			m1_ddr2_memory_status_local_init_done                : out   std_logic;                                        -- local_init_done
			m1_ddr2_memory_status_local_cal_success              : out   std_logic;                                        -- local_cal_success
			m1_ddr2_memory_status_local_cal_fail                 : out   std_logic;                                        -- local_cal_fail
			m1_ddr2_oct_rdn                                      : in    std_logic                     := 'X';             -- rdn
			m1_ddr2_oct_rup                                      : in    std_logic                     := 'X';             -- rup
			m2_ddr2_i2c_scl_export                               : out   std_logic;                                        -- export
			m2_ddr2_i2c_sda_export                               : inout std_logic                     := 'X';             -- export
			m2_ddr2_memory_mem_a                                 : out   std_logic_vector(13 downto 0);                    -- mem_a
			m2_ddr2_memory_mem_ba                                : out   std_logic_vector(2 downto 0);                     -- mem_ba
			m2_ddr2_memory_mem_ck                                : out   std_logic_vector(1 downto 0);                     -- mem_ck
			m2_ddr2_memory_mem_ck_n                              : out   std_logic_vector(1 downto 0);                     -- mem_ck_n
			m2_ddr2_memory_mem_cke                               : out   std_logic_vector(0 downto 0);                     -- mem_cke
			m2_ddr2_memory_mem_cs_n                              : out   std_logic_vector(0 downto 0);                     -- mem_cs_n
			m2_ddr2_memory_mem_dm                                : out   std_logic_vector(7 downto 0);                     -- mem_dm
			m2_ddr2_memory_mem_ras_n                             : out   std_logic_vector(0 downto 0);                     -- mem_ras_n
			m2_ddr2_memory_mem_cas_n                             : out   std_logic_vector(0 downto 0);                     -- mem_cas_n
			m2_ddr2_memory_mem_we_n                              : out   std_logic_vector(0 downto 0);                     -- mem_we_n
			m2_ddr2_memory_mem_dq                                : inout std_logic_vector(63 downto 0) := (others => 'X'); -- mem_dq
			m2_ddr2_memory_mem_dqs                               : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dqs
			m2_ddr2_memory_mem_dqs_n                             : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dqs_n
			m2_ddr2_memory_mem_odt                               : out   std_logic_vector(0 downto 0);                     -- mem_odt
			m2_ddr2_memory_dll_sharing_dll_pll_locked            : in    std_logic                     := 'X';             -- dll_pll_locked
			m2_ddr2_memory_dll_sharing_dll_delayctrl             : out   std_logic_vector(5 downto 0);                     -- dll_delayctrl
			m2_ddr2_memory_pll_sharing_pll_mem_clk               : out   std_logic;                                        -- pll_mem_clk
			m2_ddr2_memory_pll_sharing_pll_write_clk             : out   std_logic;                                        -- pll_write_clk
			m2_ddr2_memory_pll_sharing_pll_locked                : out   std_logic;                                        -- pll_locked
			m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk : out   std_logic;                                        -- pll_write_clk_pre_phy_clk
			m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk          : out   std_logic;                                        -- pll_addr_cmd_clk
			m2_ddr2_memory_pll_sharing_pll_avl_clk               : out   std_logic;                                        -- pll_avl_clk
			m2_ddr2_memory_pll_sharing_pll_config_clk            : out   std_logic;                                        -- pll_config_clk
			m2_ddr2_memory_status_local_init_done                : out   std_logic;                                        -- local_init_done
			m2_ddr2_memory_status_local_cal_success              : out   std_logic;                                        -- local_cal_success
			m2_ddr2_memory_status_local_cal_fail                 : out   std_logic;                                        -- local_cal_fail
			m2_ddr2_oct_rdn                                      : in    std_logic                     := 'X';             -- rdn
			m2_ddr2_oct_rup                                      : in    std_logic                     := 'X';             -- rup
			rst_reset_n                                          : in    std_logic                     := 'X';             -- reset_n
			sd_clk_export                                        : out   std_logic;                                        -- export
			sd_cmd_export                                        : inout std_logic                     := 'X';             -- export
			sd_dat_export                                        : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			sd_wp_n_export                                       : in    std_logic                     := 'X';             -- export
			ssdp_ssdp0                                           : out   std_logic_vector(7 downto 0);                     -- ssdp0
			ssdp_ssdp1                                           : out   std_logic_vector(7 downto 0);                     -- ssdp1
			temp_scl_export                                      : out   std_logic;                                        -- export
			temp_sda_export                                      : inout std_logic                     := 'X';             -- export
			timer_1ms_external_port_export                       : out   std_logic;                                        -- export
			timer_1us_external_port_export                       : out   std_logic;                                        -- export
			tristate_conduit_tcm_address_out                     : out   std_logic_vector(25 downto 0);                    -- tcm_address_out
			tristate_conduit_tcm_read_n_out                      : out   std_logic_vector(0 downto 0);                     -- tcm_read_n_out
			tristate_conduit_tcm_write_n_out                     : out   std_logic_vector(0 downto 0);                     -- tcm_write_n_out
			tristate_conduit_tcm_data_out                        : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			tristate_conduit_tcm_chipselect_n_out                : out   std_logic_vector(0 downto 0);                     -- tcm_chipselect_n_out
			tse_clk_clk                                          : in    std_logic                     := 'X';             -- clk
			tse_led_crs                                          : out   std_logic;                                        -- crs
			tse_led_link                                         : out   std_logic;                                        -- link
			tse_led_panel_link                                   : out   std_logic;                                        -- panel_link
			tse_led_col                                          : out   std_logic;                                        -- col
			tse_led_an                                           : out   std_logic;                                        -- an
			tse_led_char_err                                     : out   std_logic;                                        -- char_err
			tse_led_disp_err                                     : out   std_logic;                                        -- disp_err
			tse_mac_mac_misc_connection_xon_gen                  : in    std_logic                     := 'X';             -- xon_gen
			tse_mac_mac_misc_connection_xoff_gen                 : in    std_logic                     := 'X';             -- xoff_gen
			tse_mac_mac_misc_connection_magic_wakeup             : out   std_logic;                                        -- magic_wakeup
			tse_mac_mac_misc_connection_magic_sleep_n            : in    std_logic                     := 'X';             -- magic_sleep_n
			tse_mac_mac_misc_connection_ff_tx_crc_fwd            : in    std_logic                     := 'X';             -- ff_tx_crc_fwd
			tse_mac_mac_misc_connection_ff_tx_septy              : out   std_logic;                                        -- ff_tx_septy
			tse_mac_mac_misc_connection_tx_ff_uflow              : out   std_logic;                                        -- tx_ff_uflow
			tse_mac_mac_misc_connection_ff_tx_a_full             : out   std_logic;                                        -- ff_tx_a_full
			tse_mac_mac_misc_connection_ff_tx_a_empty            : out   std_logic;                                        -- ff_tx_a_empty
			tse_mac_mac_misc_connection_rx_err_stat              : out   std_logic_vector(17 downto 0);                    -- rx_err_stat
			tse_mac_mac_misc_connection_rx_frm_type              : out   std_logic_vector(3 downto 0);                     -- rx_frm_type
			tse_mac_mac_misc_connection_ff_rx_dsav               : out   std_logic;                                        -- ff_rx_dsav
			tse_mac_mac_misc_connection_ff_rx_a_full             : out   std_logic;                                        -- ff_rx_a_full
			tse_mac_mac_misc_connection_ff_rx_a_empty            : out   std_logic;                                        -- ff_rx_a_empty
			tse_mac_serdes_control_connection_export             : out   std_logic;                                        -- export
			tse_mdio_mdc                                         : out   std_logic;                                        -- mdc
			tse_mdio_mdio_in                                     : in    std_logic                     := 'X';             -- mdio_in
			tse_mdio_mdio_out                                    : out   std_logic;                                        -- mdio_out
			tse_mdio_mdio_oen                                    : out   std_logic;                                        -- mdio_oen
			tse_serial_txp                                       : out   std_logic;                                        -- txp
			tse_serial_rxp                                       : in    std_logic                     := 'X'              -- rxp
		);
	end component MebX_Qsys_Project;

	component altera_conduit_bfm is
		port (
			sig_export : out std_logic_vector(3 downto 0)   -- export
		);
	end component altera_conduit_bfm;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_conduit_bfm_0002 is
		port (
			sig_export : in std_logic_vector(0 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0002;

	component altera_conduit_bfm_0003 is
		port (
			sig_export : in std_logic_vector(1 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0003;

	component altera_conduit_bfm_0004 is
		port (
			sig_export : out std_logic_vector(0 downto 0)   -- export
		);
	end component altera_conduit_bfm_0004;

	component altera_conduit_bfm_0005 is
		port (
			sig_export : out std_logic_vector(7 downto 0)   -- export
		);
	end component altera_conduit_bfm_0005;

	component altera_conduit_bfm_0006 is
		port (
			sig_export : in std_logic_vector(7 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0006;

	component altera_conduit_bfm_0007 is
		port (
			sig_export : in std_logic_vector(12 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0007;

	component altera_conduit_bfm_0008 is
		port (
			sig_export : inout std_logic_vector(0 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0008;

	component altera_conduit_bfm_0009 is
		port (
			sig_local_init_done   : in std_logic_vector(0 downto 0) := (others => 'X'); -- local_init_done
			sig_local_cal_success : in std_logic_vector(0 downto 0) := (others => 'X'); -- local_cal_success
			sig_local_cal_fail    : in std_logic_vector(0 downto 0) := (others => 'X')  -- local_cal_fail
		);
	end component altera_conduit_bfm_0009;

	component altera_conduit_bfm_0010 is
		port (
			sig_rdn : out std_logic_vector(0 downto 0);  -- rdn
			sig_rup : out std_logic_vector(0 downto 0)   -- rup
		);
	end component altera_conduit_bfm_0010;

	component altera_conduit_bfm_0011 is
		port (
			sig_dll_pll_locked : out std_logic_vector(0 downto 0);                    -- dll_pll_locked
			sig_dll_delayctrl  : in  std_logic_vector(5 downto 0) := (others => 'X')  -- dll_delayctrl
		);
	end component altera_conduit_bfm_0011;

	component altera_conduit_bfm_0012 is
		port (
			sig_pll_mem_clk               : in std_logic_vector(0 downto 0) := (others => 'X'); -- pll_mem_clk
			sig_pll_write_clk             : in std_logic_vector(0 downto 0) := (others => 'X'); -- pll_write_clk
			sig_pll_locked                : in std_logic_vector(0 downto 0) := (others => 'X'); -- pll_locked
			sig_pll_write_clk_pre_phy_clk : in std_logic_vector(0 downto 0) := (others => 'X'); -- pll_write_clk_pre_phy_clk
			sig_pll_addr_cmd_clk          : in std_logic_vector(0 downto 0) := (others => 'X'); -- pll_addr_cmd_clk
			sig_pll_avl_clk               : in std_logic_vector(0 downto 0) := (others => 'X'); -- pll_avl_clk
			sig_pll_config_clk            : in std_logic_vector(0 downto 0) := (others => 'X')  -- pll_config_clk
		);
	end component altera_conduit_bfm_0012;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	component altera_conduit_bfm_0013 is
		port (
			sig_export : inout std_logic_vector(3 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0013;

	component altera_conduit_bfm_0014 is
		port (
			clk       : in std_logic                    := 'X';             -- clk
			reset     : in std_logic                    := 'X';             -- reset
			sig_ssdp0 : in std_logic_vector(7 downto 0) := (others => 'X'); -- ssdp0
			sig_ssdp1 : in std_logic_vector(7 downto 0) := (others => 'X')  -- ssdp1
		);
	end component altera_conduit_bfm_0014;

	component altera_conduit_bfm_0015 is
		port (
			sig_crs        : in std_logic_vector(0 downto 0) := (others => 'X'); -- crs
			sig_link       : in std_logic_vector(0 downto 0) := (others => 'X'); -- link
			sig_panel_link : in std_logic_vector(0 downto 0) := (others => 'X'); -- panel_link
			sig_col        : in std_logic_vector(0 downto 0) := (others => 'X'); -- col
			sig_an         : in std_logic_vector(0 downto 0) := (others => 'X'); -- an
			sig_char_err   : in std_logic_vector(0 downto 0) := (others => 'X'); -- char_err
			sig_disp_err   : in std_logic_vector(0 downto 0) := (others => 'X')  -- disp_err
		);
	end component altera_conduit_bfm_0015;

	component altera_conduit_bfm_0016 is
		port (
			sig_xon_gen       : out std_logic_vector(0 downto 0);                     -- xon_gen
			sig_xoff_gen      : out std_logic_vector(0 downto 0);                     -- xoff_gen
			sig_magic_wakeup  : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- magic_wakeup
			sig_magic_sleep_n : out std_logic_vector(0 downto 0);                     -- magic_sleep_n
			sig_ff_tx_crc_fwd : out std_logic_vector(0 downto 0);                     -- ff_tx_crc_fwd
			sig_ff_tx_septy   : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- ff_tx_septy
			sig_tx_ff_uflow   : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- tx_ff_uflow
			sig_ff_tx_a_full  : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- ff_tx_a_full
			sig_ff_tx_a_empty : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- ff_tx_a_empty
			sig_rx_err_stat   : in  std_logic_vector(17 downto 0) := (others => 'X'); -- rx_err_stat
			sig_rx_frm_type   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- rx_frm_type
			sig_ff_rx_dsav    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- ff_rx_dsav
			sig_ff_rx_a_full  : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- ff_rx_a_full
			sig_ff_rx_a_empty : in  std_logic_vector(0 downto 0)  := (others => 'X')  -- ff_rx_a_empty
		);
	end component altera_conduit_bfm_0016;

	component altera_conduit_bfm_0017 is
		port (
			sig_mdc      : in  std_logic_vector(0 downto 0) := (others => 'X'); -- mdc
			sig_mdio_in  : out std_logic_vector(0 downto 0);                    -- mdio_in
			sig_mdio_out : in  std_logic_vector(0 downto 0) := (others => 'X'); -- mdio_out
			sig_mdio_oen : in  std_logic_vector(0 downto 0) := (others => 'X')  -- mdio_oen
		);
	end component altera_conduit_bfm_0017;

	component altera_conduit_bfm_0018 is
		port (
			sig_txp : in  std_logic_vector(0 downto 0) := (others => 'X'); -- txp
			sig_rxp : out std_logic_vector(0 downto 0)                     -- rxp
		);
	end component altera_conduit_bfm_0018;

	component altera_external_memory_bfm_vhdl is
		generic (
			USE_CHIPSELECT           : integer := 1;
			USE_WRITE                : integer := 1;
			USE_READ                 : integer := 1;
			USE_OUTPUTENABLE         : integer := 1;
			USE_BEGINTRANSFER        : integer := 1;
			ACTIVE_LOW_BYTEENABLE    : integer := 0;
			ACTIVE_LOW_CHIPSELECT    : integer := 0;
			ACTIVE_LOW_WRITE         : integer := 0;
			ACTIVE_LOW_READ          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE  : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER : integer := 0;
			ACTIVE_LOW_RESET         : integer := 0;
			CDT_ADDRESS_W            : integer := 8;
			CDT_SYMBOL_W             : integer := 8;
			CDT_NUMSYMBOLS           : integer := 4;
			INIT_FILE                : string  := "altera_external_memory_bfm.hex";
			CDT_READ_LATENCY         : integer := 0;
			VHDL_ID                  : integer := 0
		);
		port (
			clk               : in    std_logic                     := 'X';             -- clk
			cdt_write         : in    std_logic                     := 'X';             -- tcm_write_n_out
			cdt_read          : in    std_logic                     := 'X';             -- tcm_read_n_out
			cdt_chipselect    : in    std_logic                     := 'X';             -- tcm_chipselect_n_out
			cdt_address       : in    std_logic_vector(25 downto 0) := (others => 'X'); -- tcm_address_out
			cdt_data_io       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			cdt_outputenable  : in    std_logic                     := 'X';             -- tcm_outputenable_out
			cdt_begintransfer : in    std_logic                     := 'X';             -- tcm_begintransfer_out
			cdt_byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- tcm_byteenable_out
			cdt_reset         : in    std_logic                     := 'X'              -- tcm_reset_out
		);
	end component altera_external_memory_bfm_vhdl;

	component alt_mem_if_ddr2_mem_model_top_mem_if_dm_pins_en_mem_if_dqsn_en is
		generic (
			MEM_IF_ADDR_WIDTH            : integer := 0;
			MEM_IF_ROW_ADDR_WIDTH        : integer := 0;
			MEM_IF_COL_ADDR_WIDTH        : integer := 0;
			MEM_IF_CS_PER_RANK           : integer := 0;
			MEM_IF_CONTROL_WIDTH         : integer := 0;
			MEM_IF_DQS_WIDTH             : integer := 0;
			MEM_IF_CS_WIDTH              : integer := 0;
			MEM_IF_BANKADDR_WIDTH        : integer := 0;
			MEM_IF_DQ_WIDTH              : integer := 0;
			MEM_IF_CK_WIDTH              : integer := 0;
			MEM_IF_CLK_EN_WIDTH          : integer := 0;
			MEM_TRCD                     : integer := 0;
			MEM_TRTP                     : integer := 0;
			MEM_DQS_TO_CLK_CAPTURE_DELAY : integer := 0;
			MEM_CLK_TO_DQS_CAPTURE_DELAY : integer := 0;
			MEM_IF_ODT_WIDTH             : integer := 0;
			MEM_MIRROR_ADDRESSING_DEC    : integer := 0;
			MEM_REGDIMM_ENABLED          : boolean := false;
			DEVICE_DEPTH                 : integer := 1;
			MEM_GUARANTEED_WRITE_INIT    : boolean := false;
			MEM_VERBOSE                  : boolean := true;
			MEM_INIT_EN                  : boolean := false;
			MEM_INIT_FILE                : string  := "";
			DAT_DATA_WIDTH               : integer := 32
		);
		port (
			mem_a     : in    std_logic_vector(13 downto 0) := (others => 'X'); -- mem_a
			mem_ba    : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- mem_ba
			mem_ck    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- mem_ck
			mem_ck_n  : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- mem_ck_n
			mem_cke   : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_cke
			mem_cs_n  : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_cs_n
			mem_dm    : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dm
			mem_ras_n : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_ras_n
			mem_cas_n : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_cas_n
			mem_we_n  : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_we_n
			mem_dq    : inout std_logic_vector(63 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs   : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt   : in    std_logic_vector(0 downto 0)  := (others => 'X')  -- mem_odt
		);
	end component alt_mem_if_ddr2_mem_model_top_mem_if_dm_pins_en_mem_if_dqsn_en;

	component altera_tristate_conduit_bridge_translator is
		port (
			in_tcm_address_out      : in    std_logic_vector(25 downto 0) := (others => 'X'); -- tcm_address_out
			in_tcm_read_n_out       : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tcm_read_n_out
			in_tcm_write_n_out      : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tcm_write_n_out
			in_tcm_data_out         : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			in_tcm_chipselect_n_out : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tcm_chipselect_n_out
			tcm_address_out         : out   std_logic_vector(25 downto 0);                    -- tcm_address_out
			tcm_read_n_out          : out   std_logic_vector(0 downto 0);                     -- tcm_read_n_out
			tcm_write_n_out         : out   std_logic_vector(0 downto 0);                     -- tcm_write_n_out
			tcm_data_out            : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			tcm_chipselect_n_out    : out   std_logic_vector(0 downto 0)                      -- tcm_chipselect_n_out
		);
	end component altera_tristate_conduit_bridge_translator;

	signal mebx_qsys_project_inst_clk50_bfm_clk_clk                                     : std_logic;                     -- MebX_Qsys_Project_inst_clk50_bfm:clk -> [MebX_Qsys_Project_inst:clk50_clk, MebX_Qsys_Project_inst_rst_bfm:clk, MebX_Qsys_Project_inst_ssdp_bfm:clk]
	signal ext_flash_external_mem_bfm_clk_bfm_clk_clk                                   : std_logic;                     -- ext_flash_external_mem_bfm_clk_bfm:clk -> ext_flash_external_mem_bfm:clk
	signal mebx_qsys_project_inst_m1_ddr2_memory_pll_ref_clk_bfm_clk_clk                : std_logic;                     -- MebX_Qsys_Project_inst_m1_ddr2_memory_pll_ref_clk_bfm:clk -> MebX_Qsys_Project_inst:m1_ddr2_memory_pll_ref_clk_clk
	signal mebx_qsys_project_inst_tse_clk_bfm_clk_clk                                   : std_logic;                     -- MebX_Qsys_Project_inst_tse_clk_bfm:clk -> MebX_Qsys_Project_inst:tse_clk_clk
	signal mebx_qsys_project_inst_button_bfm_conduit_export                             : std_logic_vector(3 downto 0);  -- MebX_Qsys_Project_inst_button_bfm:sig_export -> MebX_Qsys_Project_inst:button_export
	signal mebx_qsys_project_inst_csense_adc_fo_export                                  : std_logic;                     -- MebX_Qsys_Project_inst:csense_adc_fo_export -> MebX_Qsys_Project_inst_csense_adc_fo_bfm:sig_export
	signal mebx_qsys_project_inst_csense_cs_n_export                                    : std_logic_vector(1 downto 0);  -- MebX_Qsys_Project_inst:csense_cs_n_export -> MebX_Qsys_Project_inst_csense_cs_n_bfm:sig_export
	signal mebx_qsys_project_inst_csense_sck_export                                     : std_logic;                     -- MebX_Qsys_Project_inst:csense_sck_export -> MebX_Qsys_Project_inst_csense_sck_bfm:sig_export
	signal mebx_qsys_project_inst_csense_sdi_export                                     : std_logic;                     -- MebX_Qsys_Project_inst:csense_sdi_export -> MebX_Qsys_Project_inst_csense_sdi_bfm:sig_export
	signal mebx_qsys_project_inst_csense_sdo_bfm_conduit_export                         : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst_csense_sdo_bfm:sig_export -> MebX_Qsys_Project_inst:csense_sdo_export
	signal mebx_qsys_project_inst_dip_bfm_conduit_export                                : std_logic_vector(7 downto 0);  -- MebX_Qsys_Project_inst_dip_bfm:sig_export -> MebX_Qsys_Project_inst:dip_export
	signal mebx_qsys_project_inst_eth_rst_export                                        : std_logic;                     -- MebX_Qsys_Project_inst:eth_rst_export -> MebX_Qsys_Project_inst_eth_rst_bfm:sig_export
	signal mebx_qsys_project_inst_ext_bfm_conduit_export                                : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst_ext_bfm:sig_export -> MebX_Qsys_Project_inst:ext_export
	signal mebx_qsys_project_inst_led_de4_export                                        : std_logic_vector(7 downto 0);  -- MebX_Qsys_Project_inst:led_de4_export -> MebX_Qsys_Project_inst_led_de4_bfm:sig_export
	signal mebx_qsys_project_inst_led_painel_export                                     : std_logic_vector(12 downto 0); -- MebX_Qsys_Project_inst:led_painel_export -> MebX_Qsys_Project_inst_led_painel_bfm:sig_export
	signal mebx_qsys_project_inst_m1_ddr2_i2c_scl_export                                : std_logic;                     -- MebX_Qsys_Project_inst:m1_ddr2_i2c_scl_export -> MebX_Qsys_Project_inst_m1_ddr2_i2c_scl_bfm:sig_export
	signal mebx_qsys_project_inst_m1_ddr2_i2c_sda_export                                : std_logic;                     -- [] -> [MebX_Qsys_Project_inst:m1_ddr2_i2c_sda_export, MebX_Qsys_Project_inst_m1_ddr2_i2c_sda_bfm:sig_export]
	signal mebx_qsys_project_inst_m1_ddr2_memory_status_local_cal_fail                  : std_logic;                     -- MebX_Qsys_Project_inst:m1_ddr2_memory_status_local_cal_fail -> MebX_Qsys_Project_inst_m1_ddr2_memory_status_bfm:sig_local_cal_fail
	signal mebx_qsys_project_inst_m1_ddr2_memory_status_local_init_done                 : std_logic;                     -- MebX_Qsys_Project_inst:m1_ddr2_memory_status_local_init_done -> MebX_Qsys_Project_inst_m1_ddr2_memory_status_bfm:sig_local_init_done
	signal mebx_qsys_project_inst_m1_ddr2_memory_status_local_cal_success               : std_logic;                     -- MebX_Qsys_Project_inst:m1_ddr2_memory_status_local_cal_success -> MebX_Qsys_Project_inst_m1_ddr2_memory_status_bfm:sig_local_cal_success
	signal mebx_qsys_project_inst_m1_ddr2_oct_bfm_conduit_rup                           : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst_m1_ddr2_oct_bfm:sig_rup -> MebX_Qsys_Project_inst:m1_ddr2_oct_rup
	signal mebx_qsys_project_inst_m1_ddr2_oct_bfm_conduit_rdn                           : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst_m1_ddr2_oct_bfm:sig_rdn -> MebX_Qsys_Project_inst:m1_ddr2_oct_rdn
	signal mebx_qsys_project_inst_m2_ddr2_i2c_scl_export                                : std_logic;                     -- MebX_Qsys_Project_inst:m2_ddr2_i2c_scl_export -> MebX_Qsys_Project_inst_m2_ddr2_i2c_scl_bfm:sig_export
	signal mebx_qsys_project_inst_m2_ddr2_i2c_sda_export                                : std_logic;                     -- [] -> [MebX_Qsys_Project_inst:m2_ddr2_i2c_sda_export, MebX_Qsys_Project_inst_m2_ddr2_i2c_sda_bfm:sig_export]
	signal mebx_qsys_project_inst_m2_ddr2_memory_dll_sharing_bfm_conduit_dll_pll_locked : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst_m2_ddr2_memory_dll_sharing_bfm:sig_dll_pll_locked -> MebX_Qsys_Project_inst:m2_ddr2_memory_dll_sharing_dll_pll_locked
	signal mebx_qsys_project_inst_m2_ddr2_memory_dll_sharing_dll_delayctrl              : std_logic_vector(5 downto 0);  -- MebX_Qsys_Project_inst:m2_ddr2_memory_dll_sharing_dll_delayctrl -> MebX_Qsys_Project_inst_m2_ddr2_memory_dll_sharing_bfm:sig_dll_delayctrl
	signal mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_write_clk              : std_logic;                     -- MebX_Qsys_Project_inst:m2_ddr2_memory_pll_sharing_pll_write_clk -> MebX_Qsys_Project_inst_m2_ddr2_memory_pll_sharing_bfm:sig_pll_write_clk
	signal mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_avl_clk                : std_logic;                     -- MebX_Qsys_Project_inst:m2_ddr2_memory_pll_sharing_pll_avl_clk -> MebX_Qsys_Project_inst_m2_ddr2_memory_pll_sharing_bfm:sig_pll_avl_clk
	signal mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk  : std_logic;                     -- MebX_Qsys_Project_inst:m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk -> MebX_Qsys_Project_inst_m2_ddr2_memory_pll_sharing_bfm:sig_pll_write_clk_pre_phy_clk
	signal mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk           : std_logic;                     -- MebX_Qsys_Project_inst:m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk -> MebX_Qsys_Project_inst_m2_ddr2_memory_pll_sharing_bfm:sig_pll_addr_cmd_clk
	signal mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_config_clk             : std_logic;                     -- MebX_Qsys_Project_inst:m2_ddr2_memory_pll_sharing_pll_config_clk -> MebX_Qsys_Project_inst_m2_ddr2_memory_pll_sharing_bfm:sig_pll_config_clk
	signal mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_mem_clk                : std_logic;                     -- MebX_Qsys_Project_inst:m2_ddr2_memory_pll_sharing_pll_mem_clk -> MebX_Qsys_Project_inst_m2_ddr2_memory_pll_sharing_bfm:sig_pll_mem_clk
	signal mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_locked                 : std_logic;                     -- MebX_Qsys_Project_inst:m2_ddr2_memory_pll_sharing_pll_locked -> MebX_Qsys_Project_inst_m2_ddr2_memory_pll_sharing_bfm:sig_pll_locked
	signal mebx_qsys_project_inst_m2_ddr2_memory_status_local_cal_fail                  : std_logic;                     -- MebX_Qsys_Project_inst:m2_ddr2_memory_status_local_cal_fail -> MebX_Qsys_Project_inst_m2_ddr2_memory_status_bfm:sig_local_cal_fail
	signal mebx_qsys_project_inst_m2_ddr2_memory_status_local_init_done                 : std_logic;                     -- MebX_Qsys_Project_inst:m2_ddr2_memory_status_local_init_done -> MebX_Qsys_Project_inst_m2_ddr2_memory_status_bfm:sig_local_init_done
	signal mebx_qsys_project_inst_m2_ddr2_memory_status_local_cal_success               : std_logic;                     -- MebX_Qsys_Project_inst:m2_ddr2_memory_status_local_cal_success -> MebX_Qsys_Project_inst_m2_ddr2_memory_status_bfm:sig_local_cal_success
	signal mebx_qsys_project_inst_m2_ddr2_oct_bfm_conduit_rup                           : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst_m2_ddr2_oct_bfm:sig_rup -> MebX_Qsys_Project_inst:m2_ddr2_oct_rup
	signal mebx_qsys_project_inst_m2_ddr2_oct_bfm_conduit_rdn                           : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst_m2_ddr2_oct_bfm:sig_rdn -> MebX_Qsys_Project_inst:m2_ddr2_oct_rdn
	signal tristate_conduit_bridge_0_tcb_translator_out_tcm_chipselect_n_out            : std_logic_vector(0 downto 0);  -- tristate_conduit_bridge_0_tcb_translator:tcm_chipselect_n_out -> ext_flash_external_mem_bfm:cdt_chipselect
	signal tristate_conduit_bridge_0_tcb_translator_out_tcm_address_out                 : std_logic_vector(25 downto 0); -- tristate_conduit_bridge_0_tcb_translator:tcm_address_out -> ext_flash_external_mem_bfm:cdt_address
	signal ext_flash_external_mem_bfm_conduit_tcm_data_out                              : std_logic_vector(15 downto 0); -- [] -> [ext_flash_external_mem_bfm:cdt_data_io, tristate_conduit_bridge_0_tcb_translator:tcm_data_out]
	signal tristate_conduit_bridge_0_tcb_translator_out_tcm_read_n_out                  : std_logic_vector(0 downto 0);  -- tristate_conduit_bridge_0_tcb_translator:tcm_read_n_out -> ext_flash_external_mem_bfm:cdt_read
	signal tristate_conduit_bridge_0_tcb_translator_out_tcm_write_n_out                 : std_logic_vector(0 downto 0);  -- tristate_conduit_bridge_0_tcb_translator:tcm_write_n_out -> ext_flash_external_mem_bfm:cdt_write
	signal mebx_qsys_project_inst_sd_clk_export                                         : std_logic;                     -- MebX_Qsys_Project_inst:sd_clk_export -> MebX_Qsys_Project_inst_sd_clk_bfm:sig_export
	signal mebx_qsys_project_inst_sd_cmd_export                                         : std_logic;                     -- [] -> [MebX_Qsys_Project_inst:sd_cmd_export, MebX_Qsys_Project_inst_sd_cmd_bfm:sig_export]
	signal mebx_qsys_project_inst_sd_dat_export                                         : std_logic_vector(3 downto 0);  -- [] -> [MebX_Qsys_Project_inst:sd_dat_export, MebX_Qsys_Project_inst_sd_dat_bfm:sig_export]
	signal mebx_qsys_project_inst_sd_wp_n_bfm_conduit_export                            : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst_sd_wp_n_bfm:sig_export -> MebX_Qsys_Project_inst:sd_wp_n_export
	signal mebx_qsys_project_inst_ssdp_ssdp0                                            : std_logic_vector(7 downto 0);  -- MebX_Qsys_Project_inst:ssdp_ssdp0 -> MebX_Qsys_Project_inst_ssdp_bfm:sig_ssdp0
	signal mebx_qsys_project_inst_ssdp_ssdp1                                            : std_logic_vector(7 downto 0);  -- MebX_Qsys_Project_inst:ssdp_ssdp1 -> MebX_Qsys_Project_inst_ssdp_bfm:sig_ssdp1
	signal mebx_qsys_project_inst_temp_scl_export                                       : std_logic;                     -- MebX_Qsys_Project_inst:temp_scl_export -> MebX_Qsys_Project_inst_temp_scl_bfm:sig_export
	signal mebx_qsys_project_inst_temp_sda_export                                       : std_logic;                     -- [] -> [MebX_Qsys_Project_inst:temp_sda_export, MebX_Qsys_Project_inst_temp_sda_bfm:sig_export]
	signal mebx_qsys_project_inst_timer_1ms_external_port_export                        : std_logic;                     -- MebX_Qsys_Project_inst:timer_1ms_external_port_export -> MebX_Qsys_Project_inst_timer_1ms_external_port_bfm:sig_export
	signal mebx_qsys_project_inst_timer_1us_external_port_export                        : std_logic;                     -- MebX_Qsys_Project_inst:timer_1us_external_port_export -> MebX_Qsys_Project_inst_timer_1us_external_port_bfm:sig_export
	signal mebx_qsys_project_inst_tse_led_disp_err                                      : std_logic;                     -- MebX_Qsys_Project_inst:tse_led_disp_err -> MebX_Qsys_Project_inst_tse_led_bfm:sig_disp_err
	signal mebx_qsys_project_inst_tse_led_col                                           : std_logic;                     -- MebX_Qsys_Project_inst:tse_led_col -> MebX_Qsys_Project_inst_tse_led_bfm:sig_col
	signal mebx_qsys_project_inst_tse_led_crs                                           : std_logic;                     -- MebX_Qsys_Project_inst:tse_led_crs -> MebX_Qsys_Project_inst_tse_led_bfm:sig_crs
	signal mebx_qsys_project_inst_tse_led_link                                          : std_logic;                     -- MebX_Qsys_Project_inst:tse_led_link -> MebX_Qsys_Project_inst_tse_led_bfm:sig_link
	signal mebx_qsys_project_inst_tse_led_char_err                                      : std_logic;                     -- MebX_Qsys_Project_inst:tse_led_char_err -> MebX_Qsys_Project_inst_tse_led_bfm:sig_char_err
	signal mebx_qsys_project_inst_tse_led_panel_link                                    : std_logic;                     -- MebX_Qsys_Project_inst:tse_led_panel_link -> MebX_Qsys_Project_inst_tse_led_bfm:sig_panel_link
	signal mebx_qsys_project_inst_tse_led_an                                            : std_logic;                     -- MebX_Qsys_Project_inst:tse_led_an -> MebX_Qsys_Project_inst_tse_led_bfm:sig_an
	signal mebx_qsys_project_inst_tse_mac_mac_misc_connection_rx_err_stat               : std_logic_vector(17 downto 0); -- MebX_Qsys_Project_inst:tse_mac_mac_misc_connection_rx_err_stat -> MebX_Qsys_Project_inst_tse_mac_mac_misc_connection_bfm:sig_rx_err_stat
	signal mebx_qsys_project_inst_tse_mac_mac_misc_connection_rx_frm_type               : std_logic_vector(3 downto 0);  -- MebX_Qsys_Project_inst:tse_mac_mac_misc_connection_rx_frm_type -> MebX_Qsys_Project_inst_tse_mac_mac_misc_connection_bfm:sig_rx_frm_type
	signal mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_rx_a_full              : std_logic;                     -- MebX_Qsys_Project_inst:tse_mac_mac_misc_connection_ff_rx_a_full -> MebX_Qsys_Project_inst_tse_mac_mac_misc_connection_bfm:sig_ff_rx_a_full
	signal mebx_qsys_project_inst_tse_mac_mac_misc_connection_bfm_conduit_magic_sleep_n : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst_tse_mac_mac_misc_connection_bfm:sig_magic_sleep_n -> MebX_Qsys_Project_inst:tse_mac_mac_misc_connection_magic_sleep_n
	signal mebx_qsys_project_inst_tse_mac_mac_misc_connection_bfm_conduit_xoff_gen      : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst_tse_mac_mac_misc_connection_bfm:sig_xoff_gen -> MebX_Qsys_Project_inst:tse_mac_mac_misc_connection_xoff_gen
	signal mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_tx_a_full              : std_logic;                     -- MebX_Qsys_Project_inst:tse_mac_mac_misc_connection_ff_tx_a_full -> MebX_Qsys_Project_inst_tse_mac_mac_misc_connection_bfm:sig_ff_tx_a_full
	signal mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_tx_a_empty             : std_logic;                     -- MebX_Qsys_Project_inst:tse_mac_mac_misc_connection_ff_tx_a_empty -> MebX_Qsys_Project_inst_tse_mac_mac_misc_connection_bfm:sig_ff_tx_a_empty
	signal mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_rx_dsav                : std_logic;                     -- MebX_Qsys_Project_inst:tse_mac_mac_misc_connection_ff_rx_dsav -> MebX_Qsys_Project_inst_tse_mac_mac_misc_connection_bfm:sig_ff_rx_dsav
	signal mebx_qsys_project_inst_tse_mac_mac_misc_connection_magic_wakeup              : std_logic;                     -- MebX_Qsys_Project_inst:tse_mac_mac_misc_connection_magic_wakeup -> MebX_Qsys_Project_inst_tse_mac_mac_misc_connection_bfm:sig_magic_wakeup
	signal mebx_qsys_project_inst_tse_mac_mac_misc_connection_bfm_conduit_xon_gen       : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst_tse_mac_mac_misc_connection_bfm:sig_xon_gen -> MebX_Qsys_Project_inst:tse_mac_mac_misc_connection_xon_gen
	signal mebx_qsys_project_inst_tse_mac_mac_misc_connection_bfm_conduit_ff_tx_crc_fwd : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst_tse_mac_mac_misc_connection_bfm:sig_ff_tx_crc_fwd -> MebX_Qsys_Project_inst:tse_mac_mac_misc_connection_ff_tx_crc_fwd
	signal mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_tx_septy               : std_logic;                     -- MebX_Qsys_Project_inst:tse_mac_mac_misc_connection_ff_tx_septy -> MebX_Qsys_Project_inst_tse_mac_mac_misc_connection_bfm:sig_ff_tx_septy
	signal mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_rx_a_empty             : std_logic;                     -- MebX_Qsys_Project_inst:tse_mac_mac_misc_connection_ff_rx_a_empty -> MebX_Qsys_Project_inst_tse_mac_mac_misc_connection_bfm:sig_ff_rx_a_empty
	signal mebx_qsys_project_inst_tse_mac_mac_misc_connection_tx_ff_uflow               : std_logic;                     -- MebX_Qsys_Project_inst:tse_mac_mac_misc_connection_tx_ff_uflow -> MebX_Qsys_Project_inst_tse_mac_mac_misc_connection_bfm:sig_tx_ff_uflow
	signal mebx_qsys_project_inst_tse_mac_serdes_control_connection_export              : std_logic;                     -- MebX_Qsys_Project_inst:tse_mac_serdes_control_connection_export -> MebX_Qsys_Project_inst_tse_mac_serdes_control_connection_bfm:sig_export
	signal mebx_qsys_project_inst_tse_mdio_bfm_conduit_mdio_in                          : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst_tse_mdio_bfm:sig_mdio_in -> MebX_Qsys_Project_inst:tse_mdio_mdio_in
	signal mebx_qsys_project_inst_tse_mdio_mdio_oen                                     : std_logic;                     -- MebX_Qsys_Project_inst:tse_mdio_mdio_oen -> MebX_Qsys_Project_inst_tse_mdio_bfm:sig_mdio_oen
	signal mebx_qsys_project_inst_tse_mdio_mdio_out                                     : std_logic;                     -- MebX_Qsys_Project_inst:tse_mdio_mdio_out -> MebX_Qsys_Project_inst_tse_mdio_bfm:sig_mdio_out
	signal mebx_qsys_project_inst_tse_mdio_mdc                                          : std_logic;                     -- MebX_Qsys_Project_inst:tse_mdio_mdc -> MebX_Qsys_Project_inst_tse_mdio_bfm:sig_mdc
	signal mebx_qsys_project_inst_tse_serial_bfm_conduit_rxp                            : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst_tse_serial_bfm:sig_rxp -> MebX_Qsys_Project_inst:tse_serial_rxp
	signal mebx_qsys_project_inst_tse_serial_txp                                        : std_logic;                     -- MebX_Qsys_Project_inst:tse_serial_txp -> MebX_Qsys_Project_inst_tse_serial_bfm:sig_txp
	signal mebx_qsys_project_inst_tristate_conduit_tcm_chipselect_n_out                 : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:tristate_conduit_tcm_chipselect_n_out -> tristate_conduit_bridge_0_tcb_translator:in_tcm_chipselect_n_out
	signal mebx_qsys_project_inst_tristate_conduit_tcm_address_out                      : std_logic_vector(25 downto 0); -- MebX_Qsys_Project_inst:tristate_conduit_tcm_address_out -> tristate_conduit_bridge_0_tcb_translator:in_tcm_address_out
	signal mebx_qsys_project_inst_tristate_conduit_tcm_data_out                         : std_logic_vector(15 downto 0); -- [] -> [MebX_Qsys_Project_inst:tristate_conduit_tcm_data_out, tristate_conduit_bridge_0_tcb_translator:in_tcm_data_out]
	signal mebx_qsys_project_inst_tristate_conduit_tcm_read_n_out                       : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:tristate_conduit_tcm_read_n_out -> tristate_conduit_bridge_0_tcb_translator:in_tcm_read_n_out
	signal mebx_qsys_project_inst_tristate_conduit_tcm_write_n_out                      : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:tristate_conduit_tcm_write_n_out -> tristate_conduit_bridge_0_tcb_translator:in_tcm_write_n_out
	signal mebx_qsys_project_inst_m1_ddr2_memory_mem_cas_n                              : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:m1_ddr2_memory_mem_cas_n -> m1_ddr2_memory_mem_model:mem_cas_n
	signal mebx_qsys_project_inst_m1_ddr2_memory_mem_ba                                 : std_logic_vector(2 downto 0);  -- MebX_Qsys_Project_inst:m1_ddr2_memory_mem_ba -> m1_ddr2_memory_mem_model:mem_ba
	signal mebx_qsys_project_inst_m1_ddr2_memory_mem_we_n                               : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:m1_ddr2_memory_mem_we_n -> m1_ddr2_memory_mem_model:mem_we_n
	signal mebx_qsys_project_inst_m1_ddr2_memory_mem_ck                                 : std_logic_vector(1 downto 0);  -- MebX_Qsys_Project_inst:m1_ddr2_memory_mem_ck -> m1_ddr2_memory_mem_model:mem_ck
	signal mebx_qsys_project_inst_m1_ddr2_memory_mem_dm                                 : std_logic_vector(7 downto 0);  -- MebX_Qsys_Project_inst:m1_ddr2_memory_mem_dm -> m1_ddr2_memory_mem_model:mem_dm
	signal mebx_qsys_project_inst_m1_ddr2_memory_mem_dqs                                : std_logic_vector(7 downto 0);  -- [] -> [MebX_Qsys_Project_inst:m1_ddr2_memory_mem_dqs, m1_ddr2_memory_mem_model:mem_dqs]
	signal mebx_qsys_project_inst_m1_ddr2_memory_mem_dq                                 : std_logic_vector(63 downto 0); -- [] -> [MebX_Qsys_Project_inst:m1_ddr2_memory_mem_dq, m1_ddr2_memory_mem_model:mem_dq]
	signal mebx_qsys_project_inst_m1_ddr2_memory_mem_cs_n                               : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:m1_ddr2_memory_mem_cs_n -> m1_ddr2_memory_mem_model:mem_cs_n
	signal mebx_qsys_project_inst_m1_ddr2_memory_mem_a                                  : std_logic_vector(13 downto 0); -- MebX_Qsys_Project_inst:m1_ddr2_memory_mem_a -> m1_ddr2_memory_mem_model:mem_a
	signal mebx_qsys_project_inst_m1_ddr2_memory_mem_ras_n                              : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:m1_ddr2_memory_mem_ras_n -> m1_ddr2_memory_mem_model:mem_ras_n
	signal mebx_qsys_project_inst_m1_ddr2_memory_mem_dqs_n                              : std_logic_vector(7 downto 0);  -- [] -> [MebX_Qsys_Project_inst:m1_ddr2_memory_mem_dqs_n, m1_ddr2_memory_mem_model:mem_dqs_n]
	signal mebx_qsys_project_inst_m1_ddr2_memory_mem_odt                                : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:m1_ddr2_memory_mem_odt -> m1_ddr2_memory_mem_model:mem_odt
	signal mebx_qsys_project_inst_m1_ddr2_memory_mem_ck_n                               : std_logic_vector(1 downto 0);  -- MebX_Qsys_Project_inst:m1_ddr2_memory_mem_ck_n -> m1_ddr2_memory_mem_model:mem_ck_n
	signal mebx_qsys_project_inst_m1_ddr2_memory_mem_cke                                : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:m1_ddr2_memory_mem_cke -> m1_ddr2_memory_mem_model:mem_cke
	signal mebx_qsys_project_inst_m2_ddr2_memory_mem_cas_n                              : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:m2_ddr2_memory_mem_cas_n -> m2_ddr2_memory_mem_model:mem_cas_n
	signal mebx_qsys_project_inst_m2_ddr2_memory_mem_ba                                 : std_logic_vector(2 downto 0);  -- MebX_Qsys_Project_inst:m2_ddr2_memory_mem_ba -> m2_ddr2_memory_mem_model:mem_ba
	signal mebx_qsys_project_inst_m2_ddr2_memory_mem_we_n                               : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:m2_ddr2_memory_mem_we_n -> m2_ddr2_memory_mem_model:mem_we_n
	signal mebx_qsys_project_inst_m2_ddr2_memory_mem_ck                                 : std_logic_vector(1 downto 0);  -- MebX_Qsys_Project_inst:m2_ddr2_memory_mem_ck -> m2_ddr2_memory_mem_model:mem_ck
	signal mebx_qsys_project_inst_m2_ddr2_memory_mem_dm                                 : std_logic_vector(7 downto 0);  -- MebX_Qsys_Project_inst:m2_ddr2_memory_mem_dm -> m2_ddr2_memory_mem_model:mem_dm
	signal mebx_qsys_project_inst_m2_ddr2_memory_mem_dqs                                : std_logic_vector(7 downto 0);  -- [] -> [MebX_Qsys_Project_inst:m2_ddr2_memory_mem_dqs, m2_ddr2_memory_mem_model:mem_dqs]
	signal mebx_qsys_project_inst_m2_ddr2_memory_mem_dq                                 : std_logic_vector(63 downto 0); -- [] -> [MebX_Qsys_Project_inst:m2_ddr2_memory_mem_dq, m2_ddr2_memory_mem_model:mem_dq]
	signal mebx_qsys_project_inst_m2_ddr2_memory_mem_cs_n                               : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:m2_ddr2_memory_mem_cs_n -> m2_ddr2_memory_mem_model:mem_cs_n
	signal mebx_qsys_project_inst_m2_ddr2_memory_mem_a                                  : std_logic_vector(13 downto 0); -- MebX_Qsys_Project_inst:m2_ddr2_memory_mem_a -> m2_ddr2_memory_mem_model:mem_a
	signal mebx_qsys_project_inst_m2_ddr2_memory_mem_ras_n                              : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:m2_ddr2_memory_mem_ras_n -> m2_ddr2_memory_mem_model:mem_ras_n
	signal mebx_qsys_project_inst_m2_ddr2_memory_mem_dqs_n                              : std_logic_vector(7 downto 0);  -- [] -> [MebX_Qsys_Project_inst:m2_ddr2_memory_mem_dqs_n, m2_ddr2_memory_mem_model:mem_dqs_n]
	signal mebx_qsys_project_inst_m2_ddr2_memory_mem_odt                                : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:m2_ddr2_memory_mem_odt -> m2_ddr2_memory_mem_model:mem_odt
	signal mebx_qsys_project_inst_m2_ddr2_memory_mem_ck_n                               : std_logic_vector(1 downto 0);  -- MebX_Qsys_Project_inst:m2_ddr2_memory_mem_ck_n -> m2_ddr2_memory_mem_model:mem_ck_n
	signal mebx_qsys_project_inst_m2_ddr2_memory_mem_cke                                : std_logic_vector(0 downto 0);  -- MebX_Qsys_Project_inst:m2_ddr2_memory_mem_cke -> m2_ddr2_memory_mem_model:mem_cke
	signal mebx_qsys_project_inst_rst_bfm_reset_reset                                   : std_logic;                     -- MebX_Qsys_Project_inst_rst_bfm:reset -> [MebX_Qsys_Project_inst:rst_reset_n, mebx_qsys_project_inst_rst_bfm_reset_reset:in]
	signal mebx_qsys_project_inst_rst_bfm_reset_reset_ports_inv                         : std_logic;                     -- mebx_qsys_project_inst_rst_bfm_reset_reset:inv -> MebX_Qsys_Project_inst_ssdp_bfm:reset

begin

	mebx_qsys_project_inst : component MebX_Qsys_Project
		port map (
			button_export                                        => mebx_qsys_project_inst_button_bfm_conduit_export,                                --                            button.export
			clk50_clk                                            => mebx_qsys_project_inst_clk50_bfm_clk_clk,                                        --                             clk50.clk
			csense_adc_fo_export                                 => mebx_qsys_project_inst_csense_adc_fo_export,                                     --                     csense_adc_fo.export
			csense_cs_n_export                                   => mebx_qsys_project_inst_csense_cs_n_export,                                       --                       csense_cs_n.export
			csense_sck_export                                    => mebx_qsys_project_inst_csense_sck_export,                                        --                        csense_sck.export
			csense_sdi_export                                    => mebx_qsys_project_inst_csense_sdi_export,                                        --                        csense_sdi.export
			csense_sdo_export                                    => mebx_qsys_project_inst_csense_sdo_bfm_conduit_export(0),                         --                        csense_sdo.export
			dip_export                                           => mebx_qsys_project_inst_dip_bfm_conduit_export,                                   --                               dip.export
			eth_rst_export                                       => mebx_qsys_project_inst_eth_rst_export,                                           --                           eth_rst.export
			ext_export                                           => mebx_qsys_project_inst_ext_bfm_conduit_export(0),                                --                               ext.export
			led_de4_export                                       => mebx_qsys_project_inst_led_de4_export,                                           --                           led_de4.export
			led_painel_export                                    => mebx_qsys_project_inst_led_painel_export,                                        --                        led_painel.export
			m1_ddr2_i2c_scl_export                               => mebx_qsys_project_inst_m1_ddr2_i2c_scl_export,                                   --                   m1_ddr2_i2c_scl.export
			m1_ddr2_i2c_sda_export                               => mebx_qsys_project_inst_m1_ddr2_i2c_sda_export,                                   --                   m1_ddr2_i2c_sda.export
			m1_ddr2_memory_mem_a                                 => mebx_qsys_project_inst_m1_ddr2_memory_mem_a,                                     --                    m1_ddr2_memory.mem_a
			m1_ddr2_memory_mem_ba                                => mebx_qsys_project_inst_m1_ddr2_memory_mem_ba,                                    --                                  .mem_ba
			m1_ddr2_memory_mem_ck                                => mebx_qsys_project_inst_m1_ddr2_memory_mem_ck,                                    --                                  .mem_ck
			m1_ddr2_memory_mem_ck_n                              => mebx_qsys_project_inst_m1_ddr2_memory_mem_ck_n,                                  --                                  .mem_ck_n
			m1_ddr2_memory_mem_cke                               => mebx_qsys_project_inst_m1_ddr2_memory_mem_cke,                                   --                                  .mem_cke
			m1_ddr2_memory_mem_cs_n                              => mebx_qsys_project_inst_m1_ddr2_memory_mem_cs_n,                                  --                                  .mem_cs_n
			m1_ddr2_memory_mem_dm                                => mebx_qsys_project_inst_m1_ddr2_memory_mem_dm,                                    --                                  .mem_dm
			m1_ddr2_memory_mem_ras_n                             => mebx_qsys_project_inst_m1_ddr2_memory_mem_ras_n,                                 --                                  .mem_ras_n
			m1_ddr2_memory_mem_cas_n                             => mebx_qsys_project_inst_m1_ddr2_memory_mem_cas_n,                                 --                                  .mem_cas_n
			m1_ddr2_memory_mem_we_n                              => mebx_qsys_project_inst_m1_ddr2_memory_mem_we_n,                                  --                                  .mem_we_n
			m1_ddr2_memory_mem_dq                                => mebx_qsys_project_inst_m1_ddr2_memory_mem_dq,                                    --                                  .mem_dq
			m1_ddr2_memory_mem_dqs                               => mebx_qsys_project_inst_m1_ddr2_memory_mem_dqs,                                   --                                  .mem_dqs
			m1_ddr2_memory_mem_dqs_n                             => mebx_qsys_project_inst_m1_ddr2_memory_mem_dqs_n,                                 --                                  .mem_dqs_n
			m1_ddr2_memory_mem_odt                               => mebx_qsys_project_inst_m1_ddr2_memory_mem_odt,                                   --                                  .mem_odt
			m1_ddr2_memory_pll_ref_clk_clk                       => mebx_qsys_project_inst_m1_ddr2_memory_pll_ref_clk_bfm_clk_clk,                   --        m1_ddr2_memory_pll_ref_clk.clk
			m1_ddr2_memory_status_local_init_done                => mebx_qsys_project_inst_m1_ddr2_memory_status_local_init_done,                    --             m1_ddr2_memory_status.local_init_done
			m1_ddr2_memory_status_local_cal_success              => mebx_qsys_project_inst_m1_ddr2_memory_status_local_cal_success,                  --                                  .local_cal_success
			m1_ddr2_memory_status_local_cal_fail                 => mebx_qsys_project_inst_m1_ddr2_memory_status_local_cal_fail,                     --                                  .local_cal_fail
			m1_ddr2_oct_rdn                                      => mebx_qsys_project_inst_m1_ddr2_oct_bfm_conduit_rdn(0),                           --                       m1_ddr2_oct.rdn
			m1_ddr2_oct_rup                                      => mebx_qsys_project_inst_m1_ddr2_oct_bfm_conduit_rup(0),                           --                                  .rup
			m2_ddr2_i2c_scl_export                               => mebx_qsys_project_inst_m2_ddr2_i2c_scl_export,                                   --                   m2_ddr2_i2c_scl.export
			m2_ddr2_i2c_sda_export                               => mebx_qsys_project_inst_m2_ddr2_i2c_sda_export,                                   --                   m2_ddr2_i2c_sda.export
			m2_ddr2_memory_mem_a                                 => mebx_qsys_project_inst_m2_ddr2_memory_mem_a,                                     --                    m2_ddr2_memory.mem_a
			m2_ddr2_memory_mem_ba                                => mebx_qsys_project_inst_m2_ddr2_memory_mem_ba,                                    --                                  .mem_ba
			m2_ddr2_memory_mem_ck                                => mebx_qsys_project_inst_m2_ddr2_memory_mem_ck,                                    --                                  .mem_ck
			m2_ddr2_memory_mem_ck_n                              => mebx_qsys_project_inst_m2_ddr2_memory_mem_ck_n,                                  --                                  .mem_ck_n
			m2_ddr2_memory_mem_cke                               => mebx_qsys_project_inst_m2_ddr2_memory_mem_cke,                                   --                                  .mem_cke
			m2_ddr2_memory_mem_cs_n                              => mebx_qsys_project_inst_m2_ddr2_memory_mem_cs_n,                                  --                                  .mem_cs_n
			m2_ddr2_memory_mem_dm                                => mebx_qsys_project_inst_m2_ddr2_memory_mem_dm,                                    --                                  .mem_dm
			m2_ddr2_memory_mem_ras_n                             => mebx_qsys_project_inst_m2_ddr2_memory_mem_ras_n,                                 --                                  .mem_ras_n
			m2_ddr2_memory_mem_cas_n                             => mebx_qsys_project_inst_m2_ddr2_memory_mem_cas_n,                                 --                                  .mem_cas_n
			m2_ddr2_memory_mem_we_n                              => mebx_qsys_project_inst_m2_ddr2_memory_mem_we_n,                                  --                                  .mem_we_n
			m2_ddr2_memory_mem_dq                                => mebx_qsys_project_inst_m2_ddr2_memory_mem_dq,                                    --                                  .mem_dq
			m2_ddr2_memory_mem_dqs                               => mebx_qsys_project_inst_m2_ddr2_memory_mem_dqs,                                   --                                  .mem_dqs
			m2_ddr2_memory_mem_dqs_n                             => mebx_qsys_project_inst_m2_ddr2_memory_mem_dqs_n,                                 --                                  .mem_dqs_n
			m2_ddr2_memory_mem_odt                               => mebx_qsys_project_inst_m2_ddr2_memory_mem_odt,                                   --                                  .mem_odt
			m2_ddr2_memory_dll_sharing_dll_pll_locked            => mebx_qsys_project_inst_m2_ddr2_memory_dll_sharing_bfm_conduit_dll_pll_locked(0), --        m2_ddr2_memory_dll_sharing.dll_pll_locked
			m2_ddr2_memory_dll_sharing_dll_delayctrl             => mebx_qsys_project_inst_m2_ddr2_memory_dll_sharing_dll_delayctrl,                 --                                  .dll_delayctrl
			m2_ddr2_memory_pll_sharing_pll_mem_clk               => mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_mem_clk,                   --        m2_ddr2_memory_pll_sharing.pll_mem_clk
			m2_ddr2_memory_pll_sharing_pll_write_clk             => mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_write_clk,                 --                                  .pll_write_clk
			m2_ddr2_memory_pll_sharing_pll_locked                => mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_locked,                    --                                  .pll_locked
			m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk => mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk,     --                                  .pll_write_clk_pre_phy_clk
			m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk          => mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk,              --                                  .pll_addr_cmd_clk
			m2_ddr2_memory_pll_sharing_pll_avl_clk               => mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_avl_clk,                   --                                  .pll_avl_clk
			m2_ddr2_memory_pll_sharing_pll_config_clk            => mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_config_clk,                --                                  .pll_config_clk
			m2_ddr2_memory_status_local_init_done                => mebx_qsys_project_inst_m2_ddr2_memory_status_local_init_done,                    --             m2_ddr2_memory_status.local_init_done
			m2_ddr2_memory_status_local_cal_success              => mebx_qsys_project_inst_m2_ddr2_memory_status_local_cal_success,                  --                                  .local_cal_success
			m2_ddr2_memory_status_local_cal_fail                 => mebx_qsys_project_inst_m2_ddr2_memory_status_local_cal_fail,                     --                                  .local_cal_fail
			m2_ddr2_oct_rdn                                      => mebx_qsys_project_inst_m2_ddr2_oct_bfm_conduit_rdn(0),                           --                       m2_ddr2_oct.rdn
			m2_ddr2_oct_rup                                      => mebx_qsys_project_inst_m2_ddr2_oct_bfm_conduit_rup(0),                           --                                  .rup
			rst_reset_n                                          => mebx_qsys_project_inst_rst_bfm_reset_reset,                                      --                               rst.reset_n
			sd_clk_export                                        => mebx_qsys_project_inst_sd_clk_export,                                            --                            sd_clk.export
			sd_cmd_export                                        => mebx_qsys_project_inst_sd_cmd_export,                                            --                            sd_cmd.export
			sd_dat_export                                        => mebx_qsys_project_inst_sd_dat_export,                                            --                            sd_dat.export
			sd_wp_n_export                                       => mebx_qsys_project_inst_sd_wp_n_bfm_conduit_export(0),                            --                           sd_wp_n.export
			ssdp_ssdp0                                           => mebx_qsys_project_inst_ssdp_ssdp0,                                               --                              ssdp.ssdp0
			ssdp_ssdp1                                           => mebx_qsys_project_inst_ssdp_ssdp1,                                               --                                  .ssdp1
			temp_scl_export                                      => mebx_qsys_project_inst_temp_scl_export,                                          --                          temp_scl.export
			temp_sda_export                                      => mebx_qsys_project_inst_temp_sda_export,                                          --                          temp_sda.export
			timer_1ms_external_port_export                       => mebx_qsys_project_inst_timer_1ms_external_port_export,                           --           timer_1ms_external_port.export
			timer_1us_external_port_export                       => mebx_qsys_project_inst_timer_1us_external_port_export,                           --           timer_1us_external_port.export
			tristate_conduit_tcm_address_out                     => mebx_qsys_project_inst_tristate_conduit_tcm_address_out,                         --                  tristate_conduit.tcm_address_out
			tristate_conduit_tcm_read_n_out                      => mebx_qsys_project_inst_tristate_conduit_tcm_read_n_out,                          --                                  .tcm_read_n_out
			tristate_conduit_tcm_write_n_out                     => mebx_qsys_project_inst_tristate_conduit_tcm_write_n_out,                         --                                  .tcm_write_n_out
			tristate_conduit_tcm_data_out                        => mebx_qsys_project_inst_tristate_conduit_tcm_data_out,                            --                                  .tcm_data_out
			tristate_conduit_tcm_chipselect_n_out                => mebx_qsys_project_inst_tristate_conduit_tcm_chipselect_n_out,                    --                                  .tcm_chipselect_n_out
			tse_clk_clk                                          => mebx_qsys_project_inst_tse_clk_bfm_clk_clk,                                      --                           tse_clk.clk
			tse_led_crs                                          => mebx_qsys_project_inst_tse_led_crs,                                              --                           tse_led.crs
			tse_led_link                                         => mebx_qsys_project_inst_tse_led_link,                                             --                                  .link
			tse_led_panel_link                                   => mebx_qsys_project_inst_tse_led_panel_link,                                       --                                  .panel_link
			tse_led_col                                          => mebx_qsys_project_inst_tse_led_col,                                              --                                  .col
			tse_led_an                                           => mebx_qsys_project_inst_tse_led_an,                                               --                                  .an
			tse_led_char_err                                     => mebx_qsys_project_inst_tse_led_char_err,                                         --                                  .char_err
			tse_led_disp_err                                     => mebx_qsys_project_inst_tse_led_disp_err,                                         --                                  .disp_err
			tse_mac_mac_misc_connection_xon_gen                  => mebx_qsys_project_inst_tse_mac_mac_misc_connection_bfm_conduit_xon_gen(0),       --       tse_mac_mac_misc_connection.xon_gen
			tse_mac_mac_misc_connection_xoff_gen                 => mebx_qsys_project_inst_tse_mac_mac_misc_connection_bfm_conduit_xoff_gen(0),      --                                  .xoff_gen
			tse_mac_mac_misc_connection_magic_wakeup             => mebx_qsys_project_inst_tse_mac_mac_misc_connection_magic_wakeup,                 --                                  .magic_wakeup
			tse_mac_mac_misc_connection_magic_sleep_n            => mebx_qsys_project_inst_tse_mac_mac_misc_connection_bfm_conduit_magic_sleep_n(0), --                                  .magic_sleep_n
			tse_mac_mac_misc_connection_ff_tx_crc_fwd            => mebx_qsys_project_inst_tse_mac_mac_misc_connection_bfm_conduit_ff_tx_crc_fwd(0), --                                  .ff_tx_crc_fwd
			tse_mac_mac_misc_connection_ff_tx_septy              => mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_tx_septy,                  --                                  .ff_tx_septy
			tse_mac_mac_misc_connection_tx_ff_uflow              => mebx_qsys_project_inst_tse_mac_mac_misc_connection_tx_ff_uflow,                  --                                  .tx_ff_uflow
			tse_mac_mac_misc_connection_ff_tx_a_full             => mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_tx_a_full,                 --                                  .ff_tx_a_full
			tse_mac_mac_misc_connection_ff_tx_a_empty            => mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_tx_a_empty,                --                                  .ff_tx_a_empty
			tse_mac_mac_misc_connection_rx_err_stat              => mebx_qsys_project_inst_tse_mac_mac_misc_connection_rx_err_stat,                  --                                  .rx_err_stat
			tse_mac_mac_misc_connection_rx_frm_type              => mebx_qsys_project_inst_tse_mac_mac_misc_connection_rx_frm_type,                  --                                  .rx_frm_type
			tse_mac_mac_misc_connection_ff_rx_dsav               => mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_rx_dsav,                   --                                  .ff_rx_dsav
			tse_mac_mac_misc_connection_ff_rx_a_full             => mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_rx_a_full,                 --                                  .ff_rx_a_full
			tse_mac_mac_misc_connection_ff_rx_a_empty            => mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_rx_a_empty,                --                                  .ff_rx_a_empty
			tse_mac_serdes_control_connection_export             => mebx_qsys_project_inst_tse_mac_serdes_control_connection_export,                 -- tse_mac_serdes_control_connection.export
			tse_mdio_mdc                                         => mebx_qsys_project_inst_tse_mdio_mdc,                                             --                          tse_mdio.mdc
			tse_mdio_mdio_in                                     => mebx_qsys_project_inst_tse_mdio_bfm_conduit_mdio_in(0),                          --                                  .mdio_in
			tse_mdio_mdio_out                                    => mebx_qsys_project_inst_tse_mdio_mdio_out,                                        --                                  .mdio_out
			tse_mdio_mdio_oen                                    => mebx_qsys_project_inst_tse_mdio_mdio_oen,                                        --                                  .mdio_oen
			tse_serial_txp                                       => mebx_qsys_project_inst_tse_serial_txp,                                           --                        tse_serial.txp
			tse_serial_rxp                                       => mebx_qsys_project_inst_tse_serial_bfm_conduit_rxp(0)                             --                                  .rxp
		);

	mebx_qsys_project_inst_button_bfm : component altera_conduit_bfm
		port map (
			sig_export => mebx_qsys_project_inst_button_bfm_conduit_export  -- conduit.export
		);

	mebx_qsys_project_inst_clk50_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => mebx_qsys_project_inst_clk50_bfm_clk_clk  -- clk.clk
		);

	mebx_qsys_project_inst_csense_adc_fo_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export(0) => mebx_qsys_project_inst_csense_adc_fo_export  -- conduit.export
		);

	mebx_qsys_project_inst_csense_cs_n_bfm : component altera_conduit_bfm_0003
		port map (
			sig_export => mebx_qsys_project_inst_csense_cs_n_export  -- conduit.export
		);

	mebx_qsys_project_inst_csense_sck_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export(0) => mebx_qsys_project_inst_csense_sck_export  -- conduit.export
		);

	mebx_qsys_project_inst_csense_sdi_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export(0) => mebx_qsys_project_inst_csense_sdi_export  -- conduit.export
		);

	mebx_qsys_project_inst_csense_sdo_bfm : component altera_conduit_bfm_0004
		port map (
			sig_export => mebx_qsys_project_inst_csense_sdo_bfm_conduit_export  -- conduit.export
		);

	mebx_qsys_project_inst_dip_bfm : component altera_conduit_bfm_0005
		port map (
			sig_export => mebx_qsys_project_inst_dip_bfm_conduit_export  -- conduit.export
		);

	mebx_qsys_project_inst_eth_rst_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export(0) => mebx_qsys_project_inst_eth_rst_export  -- conduit.export
		);

	mebx_qsys_project_inst_ext_bfm : component altera_conduit_bfm_0004
		port map (
			sig_export => mebx_qsys_project_inst_ext_bfm_conduit_export  -- conduit.export
		);

	mebx_qsys_project_inst_led_de4_bfm : component altera_conduit_bfm_0006
		port map (
			sig_export => mebx_qsys_project_inst_led_de4_export  -- conduit.export
		);

	mebx_qsys_project_inst_led_painel_bfm : component altera_conduit_bfm_0007
		port map (
			sig_export => mebx_qsys_project_inst_led_painel_export  -- conduit.export
		);

	mebx_qsys_project_inst_m1_ddr2_i2c_scl_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export(0) => mebx_qsys_project_inst_m1_ddr2_i2c_scl_export  -- conduit.export
		);

	mebx_qsys_project_inst_m1_ddr2_i2c_sda_bfm : component altera_conduit_bfm_0008
		port map (
			sig_export(0) => mebx_qsys_project_inst_m1_ddr2_i2c_sda_export  -- conduit.export
		);

	mebx_qsys_project_inst_m1_ddr2_memory_pll_ref_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => mebx_qsys_project_inst_m1_ddr2_memory_pll_ref_clk_bfm_clk_clk  -- clk.clk
		);

	mebx_qsys_project_inst_m1_ddr2_memory_status_bfm : component altera_conduit_bfm_0009
		port map (
			sig_local_init_done(0)   => mebx_qsys_project_inst_m1_ddr2_memory_status_local_init_done,   -- conduit.local_init_done
			sig_local_cal_success(0) => mebx_qsys_project_inst_m1_ddr2_memory_status_local_cal_success, --        .local_cal_success
			sig_local_cal_fail(0)    => mebx_qsys_project_inst_m1_ddr2_memory_status_local_cal_fail     --        .local_cal_fail
		);

	mebx_qsys_project_inst_m1_ddr2_oct_bfm : component altera_conduit_bfm_0010
		port map (
			sig_rdn => mebx_qsys_project_inst_m1_ddr2_oct_bfm_conduit_rdn, -- conduit.rdn
			sig_rup => mebx_qsys_project_inst_m1_ddr2_oct_bfm_conduit_rup  --        .rup
		);

	mebx_qsys_project_inst_m2_ddr2_i2c_scl_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export(0) => mebx_qsys_project_inst_m2_ddr2_i2c_scl_export  -- conduit.export
		);

	mebx_qsys_project_inst_m2_ddr2_i2c_sda_bfm : component altera_conduit_bfm_0008
		port map (
			sig_export(0) => mebx_qsys_project_inst_m2_ddr2_i2c_sda_export  -- conduit.export
		);

	mebx_qsys_project_inst_m2_ddr2_memory_dll_sharing_bfm : component altera_conduit_bfm_0011
		port map (
			sig_dll_pll_locked => mebx_qsys_project_inst_m2_ddr2_memory_dll_sharing_bfm_conduit_dll_pll_locked, -- conduit.dll_pll_locked
			sig_dll_delayctrl  => mebx_qsys_project_inst_m2_ddr2_memory_dll_sharing_dll_delayctrl               --        .dll_delayctrl
		);

	mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_bfm : component altera_conduit_bfm_0012
		port map (
			sig_pll_mem_clk(0)               => mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_mem_clk,               -- conduit.pll_mem_clk
			sig_pll_write_clk(0)             => mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_write_clk,             --        .pll_write_clk
			sig_pll_locked(0)                => mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_locked,                --        .pll_locked
			sig_pll_write_clk_pre_phy_clk(0) => mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk, --        .pll_write_clk_pre_phy_clk
			sig_pll_addr_cmd_clk(0)          => mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk,          --        .pll_addr_cmd_clk
			sig_pll_avl_clk(0)               => mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_avl_clk,               --        .pll_avl_clk
			sig_pll_config_clk(0)            => mebx_qsys_project_inst_m2_ddr2_memory_pll_sharing_pll_config_clk             --        .pll_config_clk
		);

	mebx_qsys_project_inst_m2_ddr2_memory_status_bfm : component altera_conduit_bfm_0009
		port map (
			sig_local_init_done(0)   => mebx_qsys_project_inst_m2_ddr2_memory_status_local_init_done,   -- conduit.local_init_done
			sig_local_cal_success(0) => mebx_qsys_project_inst_m2_ddr2_memory_status_local_cal_success, --        .local_cal_success
			sig_local_cal_fail(0)    => mebx_qsys_project_inst_m2_ddr2_memory_status_local_cal_fail     --        .local_cal_fail
		);

	mebx_qsys_project_inst_m2_ddr2_oct_bfm : component altera_conduit_bfm_0010
		port map (
			sig_rdn => mebx_qsys_project_inst_m2_ddr2_oct_bfm_conduit_rdn, -- conduit.rdn
			sig_rup => mebx_qsys_project_inst_m2_ddr2_oct_bfm_conduit_rup  --        .rup
		);

	mebx_qsys_project_inst_rst_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => mebx_qsys_project_inst_rst_bfm_reset_reset, -- reset.reset_n
			clk   => mebx_qsys_project_inst_clk50_bfm_clk_clk    --   clk.clk
		);

	mebx_qsys_project_inst_sd_clk_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export(0) => mebx_qsys_project_inst_sd_clk_export  -- conduit.export
		);

	mebx_qsys_project_inst_sd_cmd_bfm : component altera_conduit_bfm_0008
		port map (
			sig_export(0) => mebx_qsys_project_inst_sd_cmd_export  -- conduit.export
		);

	mebx_qsys_project_inst_sd_dat_bfm : component altera_conduit_bfm_0013
		port map (
			sig_export => mebx_qsys_project_inst_sd_dat_export  -- conduit.export
		);

	mebx_qsys_project_inst_sd_wp_n_bfm : component altera_conduit_bfm_0004
		port map (
			sig_export => mebx_qsys_project_inst_sd_wp_n_bfm_conduit_export  -- conduit.export
		);

	mebx_qsys_project_inst_ssdp_bfm : component altera_conduit_bfm_0014
		port map (
			clk       => mebx_qsys_project_inst_clk50_bfm_clk_clk,             --     clk.clk
			reset     => mebx_qsys_project_inst_rst_bfm_reset_reset_ports_inv, --   reset.reset
			sig_ssdp0 => mebx_qsys_project_inst_ssdp_ssdp0,                    -- conduit.ssdp0
			sig_ssdp1 => mebx_qsys_project_inst_ssdp_ssdp1                     --        .ssdp1
		);

	mebx_qsys_project_inst_temp_scl_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export(0) => mebx_qsys_project_inst_temp_scl_export  -- conduit.export
		);

	mebx_qsys_project_inst_temp_sda_bfm : component altera_conduit_bfm_0008
		port map (
			sig_export(0) => mebx_qsys_project_inst_temp_sda_export  -- conduit.export
		);

	mebx_qsys_project_inst_timer_1ms_external_port_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export(0) => mebx_qsys_project_inst_timer_1ms_external_port_export  -- conduit.export
		);

	mebx_qsys_project_inst_timer_1us_external_port_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export(0) => mebx_qsys_project_inst_timer_1us_external_port_export  -- conduit.export
		);

	mebx_qsys_project_inst_tse_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => mebx_qsys_project_inst_tse_clk_bfm_clk_clk  -- clk.clk
		);

	mebx_qsys_project_inst_tse_led_bfm : component altera_conduit_bfm_0015
		port map (
			sig_crs(0)        => mebx_qsys_project_inst_tse_led_crs,        -- conduit.crs
			sig_link(0)       => mebx_qsys_project_inst_tse_led_link,       --        .link
			sig_panel_link(0) => mebx_qsys_project_inst_tse_led_panel_link, --        .panel_link
			sig_col(0)        => mebx_qsys_project_inst_tse_led_col,        --        .col
			sig_an(0)         => mebx_qsys_project_inst_tse_led_an,         --        .an
			sig_char_err(0)   => mebx_qsys_project_inst_tse_led_char_err,   --        .char_err
			sig_disp_err(0)   => mebx_qsys_project_inst_tse_led_disp_err    --        .disp_err
		);

	mebx_qsys_project_inst_tse_mac_mac_misc_connection_bfm : component altera_conduit_bfm_0016
		port map (
			sig_xon_gen          => mebx_qsys_project_inst_tse_mac_mac_misc_connection_bfm_conduit_xon_gen,       -- conduit.xon_gen
			sig_xoff_gen         => mebx_qsys_project_inst_tse_mac_mac_misc_connection_bfm_conduit_xoff_gen,      --        .xoff_gen
			sig_magic_wakeup(0)  => mebx_qsys_project_inst_tse_mac_mac_misc_connection_magic_wakeup,              --        .magic_wakeup
			sig_magic_sleep_n    => mebx_qsys_project_inst_tse_mac_mac_misc_connection_bfm_conduit_magic_sleep_n, --        .magic_sleep_n
			sig_ff_tx_crc_fwd    => mebx_qsys_project_inst_tse_mac_mac_misc_connection_bfm_conduit_ff_tx_crc_fwd, --        .ff_tx_crc_fwd
			sig_ff_tx_septy(0)   => mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_tx_septy,               --        .ff_tx_septy
			sig_tx_ff_uflow(0)   => mebx_qsys_project_inst_tse_mac_mac_misc_connection_tx_ff_uflow,               --        .tx_ff_uflow
			sig_ff_tx_a_full(0)  => mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_tx_a_full,              --        .ff_tx_a_full
			sig_ff_tx_a_empty(0) => mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_tx_a_empty,             --        .ff_tx_a_empty
			sig_rx_err_stat      => mebx_qsys_project_inst_tse_mac_mac_misc_connection_rx_err_stat,               --        .rx_err_stat
			sig_rx_frm_type      => mebx_qsys_project_inst_tse_mac_mac_misc_connection_rx_frm_type,               --        .rx_frm_type
			sig_ff_rx_dsav(0)    => mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_rx_dsav,                --        .ff_rx_dsav
			sig_ff_rx_a_full(0)  => mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_rx_a_full,              --        .ff_rx_a_full
			sig_ff_rx_a_empty(0) => mebx_qsys_project_inst_tse_mac_mac_misc_connection_ff_rx_a_empty              --        .ff_rx_a_empty
		);

	mebx_qsys_project_inst_tse_mac_serdes_control_connection_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export(0) => mebx_qsys_project_inst_tse_mac_serdes_control_connection_export  -- conduit.export
		);

	mebx_qsys_project_inst_tse_mdio_bfm : component altera_conduit_bfm_0017
		port map (
			sig_mdc(0)      => mebx_qsys_project_inst_tse_mdio_mdc,                 -- conduit.mdc
			sig_mdio_in     => mebx_qsys_project_inst_tse_mdio_bfm_conduit_mdio_in, --        .mdio_in
			sig_mdio_out(0) => mebx_qsys_project_inst_tse_mdio_mdio_out,            --        .mdio_out
			sig_mdio_oen(0) => mebx_qsys_project_inst_tse_mdio_mdio_oen             --        .mdio_oen
		);

	mebx_qsys_project_inst_tse_serial_bfm : component altera_conduit_bfm_0018
		port map (
			sig_txp(0) => mebx_qsys_project_inst_tse_serial_txp,             -- conduit.txp
			sig_rxp    => mebx_qsys_project_inst_tse_serial_bfm_conduit_rxp  --        .rxp
		);

	ext_flash_external_mem_bfm : component altera_external_memory_bfm_vhdl
		generic map (
			USE_CHIPSELECT           => 1,
			USE_WRITE                => 1,
			USE_READ                 => 1,
			USE_OUTPUTENABLE         => 0,
			USE_BEGINTRANSFER        => 0,
			ACTIVE_LOW_BYTEENABLE    => 0,
			ACTIVE_LOW_CHIPSELECT    => 1,
			ACTIVE_LOW_WRITE         => 1,
			ACTIVE_LOW_READ          => 1,
			ACTIVE_LOW_OUTPUTENABLE  => 0,
			ACTIVE_LOW_BEGINTRANSFER => 0,
			ACTIVE_LOW_RESET         => 0,
			CDT_ADDRESS_W            => 26,
			CDT_SYMBOL_W             => 8,
			CDT_NUMSYMBOLS           => 2,
			INIT_FILE                => "altera_external_memory_bfm.hex",
			CDT_READ_LATENCY         => 0,
			VHDL_ID                  => 0
		)
		port map (
			clk               => ext_flash_external_mem_bfm_clk_bfm_clk_clk,                           --     clk.clk
			cdt_write         => tristate_conduit_bridge_0_tcb_translator_out_tcm_write_n_out(0),      -- conduit.tcm_write_n_out
			cdt_read          => tristate_conduit_bridge_0_tcb_translator_out_tcm_read_n_out(0),       --        .tcm_read_n_out
			cdt_chipselect    => tristate_conduit_bridge_0_tcb_translator_out_tcm_chipselect_n_out(0), --        .tcm_chipselect_n_out
			cdt_address       => tristate_conduit_bridge_0_tcb_translator_out_tcm_address_out,         --        .tcm_address_out
			cdt_data_io       => ext_flash_external_mem_bfm_conduit_tcm_data_out,                      --        .tcm_data_out
			cdt_outputenable  => '0',                                                                  -- (terminated)
			cdt_begintransfer => '0',                                                                  -- (terminated)
			cdt_byteenable    => "11",                                                                 -- (terminated)
			cdt_reset         => '0'                                                                   -- (terminated)
		);

	ext_flash_external_mem_bfm_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 100000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => ext_flash_external_mem_bfm_clk_bfm_clk_clk  -- clk.clk
		);

	m1_ddr2_memory_mem_model : component alt_mem_if_ddr2_mem_model_top_mem_if_dm_pins_en_mem_if_dqsn_en
		generic map (
			MEM_IF_ADDR_WIDTH            => 14,
			MEM_IF_ROW_ADDR_WIDTH        => 14,
			MEM_IF_COL_ADDR_WIDTH        => 10,
			MEM_IF_CS_PER_RANK           => 1,
			MEM_IF_CONTROL_WIDTH         => 1,
			MEM_IF_DQS_WIDTH             => 8,
			MEM_IF_CS_WIDTH              => 1,
			MEM_IF_BANKADDR_WIDTH        => 3,
			MEM_IF_DQ_WIDTH              => 64,
			MEM_IF_CK_WIDTH              => 2,
			MEM_IF_CLK_EN_WIDTH          => 1,
			MEM_TRCD                     => 6,
			MEM_TRTP                     => 3,
			MEM_DQS_TO_CLK_CAPTURE_DELAY => 100,
			MEM_CLK_TO_DQS_CAPTURE_DELAY => 100000,
			MEM_IF_ODT_WIDTH             => 1,
			MEM_MIRROR_ADDRESSING_DEC    => 0,
			MEM_REGDIMM_ENABLED          => false,
			DEVICE_DEPTH                 => 1,
			MEM_GUARANTEED_WRITE_INIT    => false,
			MEM_VERBOSE                  => true,
			MEM_INIT_EN                  => false,
			MEM_INIT_FILE                => "",
			DAT_DATA_WIDTH               => 32
		)
		port map (
			mem_a     => mebx_qsys_project_inst_m1_ddr2_memory_mem_a,     -- memory.mem_a
			mem_ba    => mebx_qsys_project_inst_m1_ddr2_memory_mem_ba,    --       .mem_ba
			mem_ck    => mebx_qsys_project_inst_m1_ddr2_memory_mem_ck,    --       .mem_ck
			mem_ck_n  => mebx_qsys_project_inst_m1_ddr2_memory_mem_ck_n,  --       .mem_ck_n
			mem_cke   => mebx_qsys_project_inst_m1_ddr2_memory_mem_cke,   --       .mem_cke
			mem_cs_n  => mebx_qsys_project_inst_m1_ddr2_memory_mem_cs_n,  --       .mem_cs_n
			mem_dm    => mebx_qsys_project_inst_m1_ddr2_memory_mem_dm,    --       .mem_dm
			mem_ras_n => mebx_qsys_project_inst_m1_ddr2_memory_mem_ras_n, --       .mem_ras_n
			mem_cas_n => mebx_qsys_project_inst_m1_ddr2_memory_mem_cas_n, --       .mem_cas_n
			mem_we_n  => mebx_qsys_project_inst_m1_ddr2_memory_mem_we_n,  --       .mem_we_n
			mem_dq    => mebx_qsys_project_inst_m1_ddr2_memory_mem_dq,    --       .mem_dq
			mem_dqs   => mebx_qsys_project_inst_m1_ddr2_memory_mem_dqs,   --       .mem_dqs
			mem_dqs_n => mebx_qsys_project_inst_m1_ddr2_memory_mem_dqs_n, --       .mem_dqs_n
			mem_odt   => mebx_qsys_project_inst_m1_ddr2_memory_mem_odt    --       .mem_odt
		);

	m2_ddr2_memory_mem_model : component alt_mem_if_ddr2_mem_model_top_mem_if_dm_pins_en_mem_if_dqsn_en
		generic map (
			MEM_IF_ADDR_WIDTH            => 14,
			MEM_IF_ROW_ADDR_WIDTH        => 14,
			MEM_IF_COL_ADDR_WIDTH        => 10,
			MEM_IF_CS_PER_RANK           => 1,
			MEM_IF_CONTROL_WIDTH         => 1,
			MEM_IF_DQS_WIDTH             => 8,
			MEM_IF_CS_WIDTH              => 1,
			MEM_IF_BANKADDR_WIDTH        => 3,
			MEM_IF_DQ_WIDTH              => 64,
			MEM_IF_CK_WIDTH              => 2,
			MEM_IF_CLK_EN_WIDTH          => 1,
			MEM_TRCD                     => 6,
			MEM_TRTP                     => 3,
			MEM_DQS_TO_CLK_CAPTURE_DELAY => 100,
			MEM_CLK_TO_DQS_CAPTURE_DELAY => 100000,
			MEM_IF_ODT_WIDTH             => 1,
			MEM_MIRROR_ADDRESSING_DEC    => 0,
			MEM_REGDIMM_ENABLED          => false,
			DEVICE_DEPTH                 => 1,
			MEM_GUARANTEED_WRITE_INIT    => false,
			MEM_VERBOSE                  => true,
			MEM_INIT_EN                  => false,
			MEM_INIT_FILE                => "",
			DAT_DATA_WIDTH               => 32
		)
		port map (
			mem_a     => mebx_qsys_project_inst_m2_ddr2_memory_mem_a,     -- memory.mem_a
			mem_ba    => mebx_qsys_project_inst_m2_ddr2_memory_mem_ba,    --       .mem_ba
			mem_ck    => mebx_qsys_project_inst_m2_ddr2_memory_mem_ck,    --       .mem_ck
			mem_ck_n  => mebx_qsys_project_inst_m2_ddr2_memory_mem_ck_n,  --       .mem_ck_n
			mem_cke   => mebx_qsys_project_inst_m2_ddr2_memory_mem_cke,   --       .mem_cke
			mem_cs_n  => mebx_qsys_project_inst_m2_ddr2_memory_mem_cs_n,  --       .mem_cs_n
			mem_dm    => mebx_qsys_project_inst_m2_ddr2_memory_mem_dm,    --       .mem_dm
			mem_ras_n => mebx_qsys_project_inst_m2_ddr2_memory_mem_ras_n, --       .mem_ras_n
			mem_cas_n => mebx_qsys_project_inst_m2_ddr2_memory_mem_cas_n, --       .mem_cas_n
			mem_we_n  => mebx_qsys_project_inst_m2_ddr2_memory_mem_we_n,  --       .mem_we_n
			mem_dq    => mebx_qsys_project_inst_m2_ddr2_memory_mem_dq,    --       .mem_dq
			mem_dqs   => mebx_qsys_project_inst_m2_ddr2_memory_mem_dqs,   --       .mem_dqs
			mem_dqs_n => mebx_qsys_project_inst_m2_ddr2_memory_mem_dqs_n, --       .mem_dqs_n
			mem_odt   => mebx_qsys_project_inst_m2_ddr2_memory_mem_odt    --       .mem_odt
		);

	tristate_conduit_bridge_0_tcb_translator : component altera_tristate_conduit_bridge_translator
		port map (
			in_tcm_address_out      => mebx_qsys_project_inst_tristate_conduit_tcm_address_out,           --  in.tcm_address_out
			in_tcm_read_n_out       => mebx_qsys_project_inst_tristate_conduit_tcm_read_n_out,            --    .tcm_read_n_out
			in_tcm_write_n_out      => mebx_qsys_project_inst_tristate_conduit_tcm_write_n_out,           --    .tcm_write_n_out
			in_tcm_data_out         => mebx_qsys_project_inst_tristate_conduit_tcm_data_out,              --    .tcm_data_out
			in_tcm_chipselect_n_out => mebx_qsys_project_inst_tristate_conduit_tcm_chipselect_n_out,      --    .tcm_chipselect_n_out
			tcm_address_out         => tristate_conduit_bridge_0_tcb_translator_out_tcm_address_out,      -- out.tcm_address_out
			tcm_read_n_out          => tristate_conduit_bridge_0_tcb_translator_out_tcm_read_n_out,       --    .tcm_read_n_out
			tcm_write_n_out         => tristate_conduit_bridge_0_tcb_translator_out_tcm_write_n_out,      --    .tcm_write_n_out
			tcm_data_out            => ext_flash_external_mem_bfm_conduit_tcm_data_out,                   --    .tcm_data_out
			tcm_chipselect_n_out    => tristate_conduit_bridge_0_tcb_translator_out_tcm_chipselect_n_out  --    .tcm_chipselect_n_out
		);

	mebx_qsys_project_inst_rst_bfm_reset_reset_ports_inv <= not mebx_qsys_project_inst_rst_bfm_reset_reset;

end architecture rtl; -- of MebX_Qsys_Project_tb
