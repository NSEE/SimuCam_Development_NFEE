LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.ALL;

ENTITY SEVEN_SEG_REGISTER IS
	PORT (
		CLK : IN STD_LOGIC;
		RST : IN STD_LOGIC;
		
		DATA_IN_AVALON : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		ADDRESS_IN_AVALON : IN  STD_LOGIC;
		ENABLE_DATA_IN_AVALON : IN  STD_LOGIC;
		
		SEG_DATA    : OUT UNSIGNED(7 DOWNTO 0);
		SEG1_ON_OFF : OUT STD_LOGIC;
		SEG1_UPDATE : OUT STD_LOGIC;
		SEG1_TEST   : OUT STD_LOGIC;
		SEG0_ON_OFF : OUT STD_LOGIC;
		SEG0_UPDATE : OUT STD_LOGIC;
		SEG0_TEST   : OUT STD_LOGIC

	);
END SEVEN_SEG_REGISTER;

ARCHITECTURE BEHAVIOUR OF SEVEN_SEG_REGISTER IS

	TYPE REG_SSDP_TYPE IS ARRAY (0 TO 1) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REG_SSDP : REG_SSDP_TYPE;

BEGIN

	GLOBAL : PROCESS(CLK, RST)
	BEGIN
	
		IF (RST = '1') THEN
			REG_SSDP(0) <= X"00_00_00_00"; -- CONTROL REGISTER
			--------------------------------------------------
			-- RESERVED | RESERVED | RESERVED | CONTROL REG --
			--------------------------------------------------
			-- CONTROL REG:
			-- 0 -> SEVEN SEGMENT DISPLAY 0 ON/OFF
			-- 1 -> SEVEN SEGMENT DISPLAY 0 UPDATE
			-- 2 -> SEVEN SEGMENT DISPLAY 0 TEST
			-- 3 -> RESERVED
			-- 4 -> SEVEN SEGMENT DISPLAY 1 ON/OFF
			-- 5 -> SEVEN SEGMENT DISPLAY 1 UPDATE
			-- 6 -> SEVEN SEGMENT DISPLAY 1 TEST
			-- 7 -> RESERVED
			REG_SSDP(1) <= X"00_00_00_00"; -- DATA REGISTER
			--------------------------------------------------
			-- RESERVED | RESERVED | RESERVED | DATA REG --
			--------------------------------------------------
			
		ELSIF (RISING_EDGE(CLK)) THEN
			IF (ENABLE_DATA_IN_AVALON = '1') THEN
				IF (ADDRESS_IN_AVALON = '0') THEN
			    	REG_SSDP(0) <= DATA_IN_AVALON;
			    ELSE
			    	REG_SSDP(1) <= DATA_IN_AVALON;
			    END IF;
				--REG_SSDP(TO_INTEGER(UNSIGNED(ADDRESS_IN_AVALON))) <= DATA_IN_AVALON;
			END IF;
		END IF;
	END PROCESS;
	
	SEG1_TEST   <= REG_SSDP(0)(6);
	SEG1_UPDATE <= REG_SSDP(0)(5);
	SEG1_ON_OFF <= REG_SSDP(0)(4);
	SEG0_TEST   <= REG_SSDP(0)(2);
	SEG0_UPDATE <= REG_SSDP(0)(1);
	SEG0_ON_OFF <= REG_SSDP(0)(0);
	SEG_DATA <= UNSIGNED(REG_SSDP(1)(7 DOWNTO 0));

END ARCHITECTURE BEHAVIOUR;

