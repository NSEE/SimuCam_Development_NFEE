package rmap_target_read_reply_header_header_crc_pkg is
	
end package rmap_target_read_reply_header_header_crc_pkg;

package body rmap_target_read_reply_header_header_crc_pkg is
	
end package body rmap_target_read_reply_header_header_crc_pkg;
