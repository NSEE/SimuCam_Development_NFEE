package rmap_memory_pkg is
	
end package rmap_memory_pkg;

package body rmap_memory_pkg is
	
end package body rmap_memory_pkg;
