-- MebX_Qsys_Project.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity MebX_Qsys_Project is
	port (
		button_export                                               : in    std_logic_vector(3 downto 0)  := (others => '0'); --                               button.export
		clk50_clk                                                   : in    std_logic                     := '0';             --                                clk50.clk
		comm_a_conduit_end_data_in_signal                           : in    std_logic                     := '0';             --                   comm_a_conduit_end.data_in_signal
		comm_a_conduit_end_data_out_signal                          : out   std_logic;                                        --                                     .data_out_signal
		comm_a_conduit_end_strobe_in_signal                         : in    std_logic                     := '0';             --                                     .strobe_in_signal
		comm_a_conduit_end_strobe_out_signal                        : out   std_logic;                                        --                                     .strobe_out_signal
		comm_a_measurements_conduit_end_measurements_channel_signal : out   std_logic_vector(7 downto 0);                     --      comm_a_measurements_conduit_end.measurements_channel_signal
		comm_a_sync_end_sync_channel_signal                         : in    std_logic                     := '0';             --                      comm_a_sync_end.sync_channel_signal
		comm_b_conduit_end_data_in_signal                           : in    std_logic                     := '0';             --                   comm_b_conduit_end.data_in_signal
		comm_b_conduit_end_data_out_signal                          : out   std_logic;                                        --                                     .data_out_signal
		comm_b_conduit_end_strobe_in_signal                         : in    std_logic                     := '0';             --                                     .strobe_in_signal
		comm_b_conduit_end_strobe_out_signal                        : out   std_logic;                                        --                                     .strobe_out_signal
		comm_b_measurements_conduit_end_measurements_channel_signal : out   std_logic_vector(7 downto 0);                     --      comm_b_measurements_conduit_end.measurements_channel_signal
		comm_b_sync_end_sync_channel_signal                         : in    std_logic                     := '0';             --                      comm_b_sync_end.sync_channel_signal
		comm_c_conduit_end_data_in_signal                           : in    std_logic                     := '0';             --                   comm_c_conduit_end.data_in_signal
		comm_c_conduit_end_data_out_signal                          : out   std_logic;                                        --                                     .data_out_signal
		comm_c_conduit_end_strobe_in_signal                         : in    std_logic                     := '0';             --                                     .strobe_in_signal
		comm_c_conduit_end_strobe_out_signal                        : out   std_logic;                                        --                                     .strobe_out_signal
		comm_c_measurements_conduit_end_measurements_channel_signal : out   std_logic_vector(7 downto 0);                     --      comm_c_measurements_conduit_end.measurements_channel_signal
		comm_c_sync_end_sync_channel_signal                         : in    std_logic                     := '0';             --                      comm_c_sync_end.sync_channel_signal
		comm_d_conduit_end_data_in_signal                           : in    std_logic                     := '0';             --                   comm_d_conduit_end.data_in_signal
		comm_d_conduit_end_data_out_signal                          : out   std_logic;                                        --                                     .data_out_signal
		comm_d_conduit_end_strobe_in_signal                         : in    std_logic                     := '0';             --                                     .strobe_in_signal
		comm_d_conduit_end_strobe_out_signal                        : out   std_logic;                                        --                                     .strobe_out_signal
		comm_d_measurements_conduit_end_measurements_channel_signal : out   std_logic_vector(7 downto 0);                     --      comm_d_measurements_conduit_end.measurements_channel_signal
		comm_d_sync_end_sync_channel_signal                         : in    std_logic                     := '0';             --                      comm_d_sync_end.sync_channel_signal
		comm_e_conduit_end_data_in_signal                           : in    std_logic                     := '0';             --                   comm_e_conduit_end.data_in_signal
		comm_e_conduit_end_data_out_signal                          : out   std_logic;                                        --                                     .data_out_signal
		comm_e_conduit_end_strobe_in_signal                         : in    std_logic                     := '0';             --                                     .strobe_in_signal
		comm_e_conduit_end_strobe_out_signal                        : out   std_logic;                                        --                                     .strobe_out_signal
		comm_e_measurements_conduit_end_measurements_channel_signal : out   std_logic_vector(7 downto 0);                     --      comm_e_measurements_conduit_end.measurements_channel_signal
		comm_e_sync_end_sync_channel_signal                         : in    std_logic                     := '0';             --                      comm_e_sync_end.sync_channel_signal
		comm_f_conduit_end_data_in_signal                           : in    std_logic                     := '0';             --                   comm_f_conduit_end.data_in_signal
		comm_f_conduit_end_data_out_signal                          : out   std_logic;                                        --                                     .data_out_signal
		comm_f_conduit_end_strobe_in_signal                         : in    std_logic                     := '0';             --                                     .strobe_in_signal
		comm_f_conduit_end_strobe_out_signal                        : out   std_logic;                                        --                                     .strobe_out_signal
		comm_f_measurements_conduit_end_measurements_channel_signal : out   std_logic_vector(7 downto 0);                     --      comm_f_measurements_conduit_end.measurements_channel_signal
		comm_f_sync_end_sync_channel_signal                         : in    std_logic                     := '0';             --                      comm_f_sync_end.sync_channel_signal
		csense_adc_fo_export                                        : out   std_logic;                                        --                        csense_adc_fo.export
		csense_cs_n_export                                          : out   std_logic_vector(1 downto 0);                     --                          csense_cs_n.export
		csense_sck_export                                           : out   std_logic;                                        --                           csense_sck.export
		csense_sdi_export                                           : out   std_logic;                                        --                           csense_sdi.export
		csense_sdo_export                                           : in    std_logic                     := '0';             --                           csense_sdo.export
		ctrl_io_lvds_export                                         : out   std_logic_vector(3 downto 0);                     --                         ctrl_io_lvds.export
		dip_export                                                  : in    std_logic_vector(7 downto 0)  := (others => '0'); --                                  dip.export
		ext_export                                                  : in    std_logic                     := '0';             --                                  ext.export
		ftdi_clk_clk                                                : in    std_logic                     := '0';             --                             ftdi_clk.clk
		led_de4_export                                              : out   std_logic_vector(7 downto 0);                     --                              led_de4.export
		led_painel_export                                           : out   std_logic_vector(20 downto 0);                    --                           led_painel.export
		m1_ddr2_i2c_scl_export                                      : out   std_logic;                                        --                      m1_ddr2_i2c_scl.export
		m1_ddr2_i2c_sda_export                                      : inout std_logic                     := '0';             --                      m1_ddr2_i2c_sda.export
		m1_ddr2_memory_mem_a                                        : out   std_logic_vector(13 downto 0);                    --                       m1_ddr2_memory.mem_a
		m1_ddr2_memory_mem_ba                                       : out   std_logic_vector(2 downto 0);                     --                                     .mem_ba
		m1_ddr2_memory_mem_ck                                       : out   std_logic_vector(1 downto 0);                     --                                     .mem_ck
		m1_ddr2_memory_mem_ck_n                                     : out   std_logic_vector(1 downto 0);                     --                                     .mem_ck_n
		m1_ddr2_memory_mem_cke                                      : out   std_logic_vector(1 downto 0);                     --                                     .mem_cke
		m1_ddr2_memory_mem_cs_n                                     : out   std_logic_vector(1 downto 0);                     --                                     .mem_cs_n
		m1_ddr2_memory_mem_dm                                       : out   std_logic_vector(7 downto 0);                     --                                     .mem_dm
		m1_ddr2_memory_mem_ras_n                                    : out   std_logic_vector(0 downto 0);                     --                                     .mem_ras_n
		m1_ddr2_memory_mem_cas_n                                    : out   std_logic_vector(0 downto 0);                     --                                     .mem_cas_n
		m1_ddr2_memory_mem_we_n                                     : out   std_logic_vector(0 downto 0);                     --                                     .mem_we_n
		m1_ddr2_memory_mem_dq                                       : inout std_logic_vector(63 downto 0) := (others => '0'); --                                     .mem_dq
		m1_ddr2_memory_mem_dqs                                      : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                     .mem_dqs
		m1_ddr2_memory_mem_dqs_n                                    : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                     .mem_dqs_n
		m1_ddr2_memory_mem_odt                                      : out   std_logic_vector(1 downto 0);                     --                                     .mem_odt
		m1_ddr2_memory_pll_ref_clk_clk                              : in    std_logic                     := '0';             --           m1_ddr2_memory_pll_ref_clk.clk
		m1_ddr2_memory_status_local_init_done                       : out   std_logic;                                        --                m1_ddr2_memory_status.local_init_done
		m1_ddr2_memory_status_local_cal_success                     : out   std_logic;                                        --                                     .local_cal_success
		m1_ddr2_memory_status_local_cal_fail                        : out   std_logic;                                        --                                     .local_cal_fail
		m1_ddr2_oct_rdn                                             : in    std_logic                     := '0';             --                          m1_ddr2_oct.rdn
		m1_ddr2_oct_rup                                             : in    std_logic                     := '0';             --                                     .rup
		m2_ddr2_i2c_scl_export                                      : out   std_logic;                                        --                      m2_ddr2_i2c_scl.export
		m2_ddr2_i2c_sda_export                                      : inout std_logic                     := '0';             --                      m2_ddr2_i2c_sda.export
		m2_ddr2_memory_mem_a                                        : out   std_logic_vector(13 downto 0);                    --                       m2_ddr2_memory.mem_a
		m2_ddr2_memory_mem_ba                                       : out   std_logic_vector(2 downto 0);                     --                                     .mem_ba
		m2_ddr2_memory_mem_ck                                       : out   std_logic_vector(1 downto 0);                     --                                     .mem_ck
		m2_ddr2_memory_mem_ck_n                                     : out   std_logic_vector(1 downto 0);                     --                                     .mem_ck_n
		m2_ddr2_memory_mem_cke                                      : out   std_logic_vector(1 downto 0);                     --                                     .mem_cke
		m2_ddr2_memory_mem_cs_n                                     : out   std_logic_vector(1 downto 0);                     --                                     .mem_cs_n
		m2_ddr2_memory_mem_dm                                       : out   std_logic_vector(7 downto 0);                     --                                     .mem_dm
		m2_ddr2_memory_mem_ras_n                                    : out   std_logic_vector(0 downto 0);                     --                                     .mem_ras_n
		m2_ddr2_memory_mem_cas_n                                    : out   std_logic_vector(0 downto 0);                     --                                     .mem_cas_n
		m2_ddr2_memory_mem_we_n                                     : out   std_logic_vector(0 downto 0);                     --                                     .mem_we_n
		m2_ddr2_memory_mem_dq                                       : inout std_logic_vector(63 downto 0) := (others => '0'); --                                     .mem_dq
		m2_ddr2_memory_mem_dqs                                      : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                     .mem_dqs
		m2_ddr2_memory_mem_dqs_n                                    : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                     .mem_dqs_n
		m2_ddr2_memory_mem_odt                                      : out   std_logic_vector(1 downto 0);                     --                                     .mem_odt
		m2_ddr2_memory_dll_sharing_dll_pll_locked                   : in    std_logic                     := '0';             --           m2_ddr2_memory_dll_sharing.dll_pll_locked
		m2_ddr2_memory_dll_sharing_dll_delayctrl                    : out   std_logic_vector(5 downto 0);                     --                                     .dll_delayctrl
		m2_ddr2_memory_pll_sharing_pll_mem_clk                      : out   std_logic;                                        --           m2_ddr2_memory_pll_sharing.pll_mem_clk
		m2_ddr2_memory_pll_sharing_pll_write_clk                    : out   std_logic;                                        --                                     .pll_write_clk
		m2_ddr2_memory_pll_sharing_pll_locked                       : out   std_logic;                                        --                                     .pll_locked
		m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk        : out   std_logic;                                        --                                     .pll_write_clk_pre_phy_clk
		m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk                 : out   std_logic;                                        --                                     .pll_addr_cmd_clk
		m2_ddr2_memory_pll_sharing_pll_avl_clk                      : out   std_logic;                                        --                                     .pll_avl_clk
		m2_ddr2_memory_pll_sharing_pll_config_clk                   : out   std_logic;                                        --                                     .pll_config_clk
		m2_ddr2_memory_status_local_init_done                       : out   std_logic;                                        --                m2_ddr2_memory_status.local_init_done
		m2_ddr2_memory_status_local_cal_success                     : out   std_logic;                                        --                                     .local_cal_success
		m2_ddr2_memory_status_local_cal_fail                        : out   std_logic;                                        --                                     .local_cal_fail
		m2_ddr2_oct_rdn                                             : in    std_logic                     := '0';             --                          m2_ddr2_oct.rdn
		m2_ddr2_oct_rup                                             : in    std_logic                     := '0';             --                                     .rup
		rs232_uart_rxd                                              : in    std_logic                     := '0';             --                           rs232_uart.rxd
		rs232_uart_txd                                              : out   std_logic;                                        --                                     .txd
		rst_reset_n                                                 : in    std_logic                     := '0';             --                                  rst.reset_n
		rst_controller_conduit_reset_input_t_reset_input_signal     : in    std_logic                     := '0';             --   rst_controller_conduit_reset_input.t_reset_input_signal
		rst_controller_conduit_simucam_reset_t_simucam_reset_signal : out   std_logic;                                        -- rst_controller_conduit_simucam_reset.t_simucam_reset_signal
		rtcc_alarm_export                                           : in    std_logic                     := '0';             --                           rtcc_alarm.export
		rtcc_cs_n_export                                            : out   std_logic;                                        --                            rtcc_cs_n.export
		rtcc_sck_export                                             : out   std_logic;                                        --                             rtcc_sck.export
		rtcc_sdi_export                                             : out   std_logic;                                        --                             rtcc_sdi.export
		rtcc_sdo_export                                             : in    std_logic                     := '0';             --                             rtcc_sdo.export
		sd_card_ip_b_SD_cmd                                         : inout std_logic                     := '0';             --                           sd_card_ip.b_SD_cmd
		sd_card_ip_b_SD_dat                                         : inout std_logic                     := '0';             --                                     .b_SD_dat
		sd_card_ip_b_SD_dat3                                        : inout std_logic                     := '0';             --                                     .b_SD_dat3
		sd_card_ip_o_SD_clock                                       : out   std_logic;                                        --                                     .o_SD_clock
		sd_card_wp_n_io_export                                      : in    std_logic                     := '0';             --                      sd_card_wp_n_io.export
		ssdp_ssdp0                                                  : out   std_logic_vector(7 downto 0);                     --                                 ssdp.ssdp0
		ssdp_ssdp1                                                  : out   std_logic_vector(7 downto 0);                     --                                     .ssdp1
		sync_in_conduit                                             : in    std_logic                     := '0';             --                              sync_in.conduit
		sync_out_conduit                                            : out   std_logic;                                        --                             sync_out.conduit
		sync_spw1_conduit                                           : out   std_logic;                                        --                            sync_spw1.conduit
		sync_spw2_conduit                                           : out   std_logic;                                        --                            sync_spw2.conduit
		sync_spw3_conduit                                           : out   std_logic;                                        --                            sync_spw3.conduit
		sync_spw4_conduit                                           : out   std_logic;                                        --                            sync_spw4.conduit
		sync_spw5_conduit                                           : out   std_logic;                                        --                            sync_spw5.conduit
		sync_spw6_conduit                                           : out   std_logic;                                        --                            sync_spw6.conduit
		sync_spw7_conduit                                           : out   std_logic;                                        --                            sync_spw7.conduit
		sync_spw8_conduit                                           : out   std_logic;                                        --                            sync_spw8.conduit
		temp_scl_export                                             : out   std_logic;                                        --                             temp_scl.export
		temp_sda_export                                             : inout std_logic                     := '0';             --                             temp_sda.export
		timer_1ms_external_port_export                              : out   std_logic;                                        --              timer_1ms_external_port.export
		timer_1us_external_port_export                              : out   std_logic;                                        --              timer_1us_external_port.export
		tristate_conduit_tcm_address_out                            : out   std_logic_vector(25 downto 0);                    --                     tristate_conduit.tcm_address_out
		tristate_conduit_tcm_read_n_out                             : out   std_logic_vector(0 downto 0);                     --                                     .tcm_read_n_out
		tristate_conduit_tcm_write_n_out                            : out   std_logic_vector(0 downto 0);                     --                                     .tcm_write_n_out
		tristate_conduit_tcm_data_out                               : inout std_logic_vector(15 downto 0) := (others => '0'); --                                     .tcm_data_out
		tristate_conduit_tcm_chipselect_n_out                       : out   std_logic_vector(0 downto 0);                     --                                     .tcm_chipselect_n_out
		umft601a_pins_umft_data_signal                              : inout std_logic_vector(31 downto 0) := (others => '0'); --                        umft601a_pins.umft_data_signal
		umft601a_pins_umft_reset_n_signal                           : out   std_logic;                                        --                                     .umft_reset_n_signal
		umft601a_pins_umft_rxf_n_signal                             : in    std_logic                     := '0';             --                                     .umft_rxf_n_signal
		umft601a_pins_umft_clock_signal                             : in    std_logic                     := '0';             --                                     .umft_clock_signal
		umft601a_pins_umft_wakeup_n_signal                          : inout std_logic                     := '0';             --                                     .umft_wakeup_n_signal
		umft601a_pins_umft_be_signal                                : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                     .umft_be_signal
		umft601a_pins_umft_txe_n_signal                             : in    std_logic                     := '0';             --                                     .umft_txe_n_signal
		umft601a_pins_umft_gpio_bus_signal                          : inout std_logic_vector(1 downto 0)  := (others => '0'); --                                     .umft_gpio_bus_signal
		umft601a_pins_umft_wr_n_signal                              : out   std_logic;                                        --                                     .umft_wr_n_signal
		umft601a_pins_umft_rd_n_signal                              : out   std_logic;                                        --                                     .umft_rd_n_signal
		umft601a_pins_umft_oe_n_signal                              : out   std_logic;                                        --                                     .umft_oe_n_signal
		umft601a_pins_umft_siwu_n_signal                            : out   std_logic                                         --                                     .umft_siwu_n_signal
	);
end entity MebX_Qsys_Project;

architecture rtl of MebX_Qsys_Project is
	component Altera_UP_SD_Card_Avalon_Interface is
		port (
			i_avalon_chip_select : in    std_logic                     := 'X';             -- chipselect
			i_avalon_address     : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			i_avalon_read        : in    std_logic                     := 'X';             -- read
			i_avalon_write       : in    std_logic                     := 'X';             -- write
			i_avalon_byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			i_avalon_writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			o_avalon_readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			o_avalon_waitrequest : out   std_logic;                                        -- waitrequest
			i_clock              : in    std_logic                     := 'X';             -- clk
			i_reset_n            : in    std_logic                     := 'X';             -- reset_n
			b_SD_cmd             : inout std_logic                     := 'X';             -- export
			b_SD_dat             : inout std_logic                     := 'X';             -- export
			b_SD_dat3            : inout std_logic                     := 'X';             -- export
			o_SD_clock           : out   std_logic                                         -- export
		);
	end component Altera_UP_SD_Card_Avalon_Interface;

	component comm_v1_80_top is
		port (
			reset_sink_reset                   : in  std_logic                      := 'X';             -- reset
			data_in                            : in  std_logic                      := 'X';             -- data_in_signal
			data_out                           : out std_logic;                                         -- data_out_signal
			strobe_in                          : in  std_logic                      := 'X';             -- strobe_in_signal
			strobe_out                         : out std_logic;                                         -- strobe_out_signal
			sync_channel                       : in  std_logic                      := 'X';             -- sync_channel_signal
			rmap_interrupt_sender_irq          : out std_logic;                                         -- irq
			buffers_interrupt_sender_irq       : out std_logic;                                         -- irq
			clock_sink_100_clk                 : in  std_logic                      := 'X';             -- clk
			clock_sink_200_clk                 : in  std_logic                      := 'X';             -- clk
			avalon_slave_windowing_address     : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- address
			avalon_slave_windowing_write       : in  std_logic                      := 'X';             -- write
			avalon_slave_windowing_read        : in  std_logic                      := 'X';             -- read
			avalon_slave_windowing_writedata   : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			avalon_slave_windowing_byteenable  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			avalon_slave_windowing_readdata    : out std_logic_vector(31 downto 0);                     -- readdata
			avalon_slave_windowing_waitrequest : out std_logic;                                         -- waitrequest
			avalon_slave_L_buffer_address      : in  std_logic_vector(20 downto 0)  := (others => 'X'); -- address
			avalon_slave_L_buffer_waitrequest  : out std_logic;                                         -- waitrequest
			avalon_slave_L_buffer_write        : in  std_logic                      := 'X';             -- write
			avalon_slave_L_buffer_writedata    : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			avalon_slave_R_buffer_address      : in  std_logic_vector(20 downto 0)  := (others => 'X'); -- address
			avalon_slave_R_buffer_write        : in  std_logic                      := 'X';             -- write
			avalon_slave_R_buffer_writedata    : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			avalon_slave_R_buffer_waitrequest  : out std_logic;                                         -- waitrequest
			measurements_channel               : out std_logic_vector(7 downto 0);                      -- measurements_channel_signal
			fee_codec_rmap_wr_waitrequest_i    : in  std_logic                      := 'X';             -- wr_waitrequest_signal
			fee_codec_rmap_readdata_i          : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata_signal
			fee_codec_rmap_rd_waitrequest_i    : in  std_logic                      := 'X';             -- rd_waitrequest_signal
			fee_codec_rmap_wr_address_o        : out std_logic_vector(31 downto 0);                     -- wr_address_signal
			fee_codec_rmap_write_o             : out std_logic;                                         -- write_signal
			fee_codec_rmap_writedata_o         : out std_logic_vector(7 downto 0);                      -- writedata_signal
			fee_codec_rmap_rd_address_o        : out std_logic_vector(31 downto 0);                     -- rd_address_signal
			fee_codec_rmap_read_o              : out std_logic;                                         -- read_signal
			fee_hk_rmap_wr_waitrequest_i       : in  std_logic                      := 'X';             -- wr_waitrequest_signal
			fee_hk_rmap_readdata_i             : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata_signal
			fee_hk_rmap_rd_waitrequest_i       : in  std_logic                      := 'X';             -- rd_waitrequest_signal
			fee_hk_rmap_wr_address_o           : out std_logic_vector(31 downto 0);                     -- wr_address_signal
			fee_hk_rmap_write_o                : out std_logic;                                         -- write_signal
			fee_hk_rmap_writedata_o            : out std_logic_vector(7 downto 0);                      -- writedata_signal
			fee_hk_rmap_rd_address_o           : out std_logic_vector(31 downto 0);                     -- rd_address_signal
			fee_hk_rmap_read_o                 : out std_logic;                                         -- read_signal
			channel_hk_timecode_control_o      : out std_logic_vector(1 downto 0);                      -- timecode_control_signal
			channel_hk_timecode_time_o         : out std_logic_vector(5 downto 0);                      -- timecode_time_signal
			channel_hk_rmap_target_status_o    : out std_logic_vector(7 downto 0);                      -- rmap_target_status_signal
			channel_hk_rmap_target_indicate_o  : out std_logic;                                         -- rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_o   : out std_logic;                                         -- spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_o   : out std_logic;                                         -- spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_o   : out std_logic;                                         -- spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_o   : out std_logic;                                         -- spw_link_disconnect_signal
			channel_hk_spw_link_running_o      : out std_logic;                                         -- spw_link_running_signal
			channel_hk_frame_counter_o         : out std_logic_vector(15 downto 0);                     -- frame_counter_signal
			channel_hk_frame_number_o          : out std_logic_vector(1 downto 0);                      -- frame_number_signal
			channel_win_mem_addr_offset_o      : out std_logic_vector(63 downto 0)                      -- win_mem_addr_offset_signal
		);
	end component comm_v1_80_top;

	component ftdi_usb3_top is
		port (
			clock_sink_clk                  : in    std_logic                      := 'X';             -- clk
			ftdi_clock_sink_clk             : in    std_logic                      := 'X';             -- clk
			reset_sink_reset                : in    std_logic                      := 'X';             -- reset
			umft_data_bus                   : inout std_logic_vector(31 downto 0)  := (others => 'X'); -- umft_data_signal
			umft_reset_n_pin                : out   std_logic;                                         -- umft_reset_n_signal
			umft_rxf_n_pin                  : in    std_logic                      := 'X';             -- umft_rxf_n_signal
			umft_clock_pin                  : in    std_logic                      := 'X';             -- umft_clock_signal
			umft_wakeup_n_pin               : inout std_logic                      := 'X';             -- umft_wakeup_n_signal
			umft_be_bus                     : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- umft_be_signal
			umft_txe_n_pin                  : in    std_logic                      := 'X';             -- umft_txe_n_signal
			umft_gpio_bus                   : inout std_logic_vector(1 downto 0)   := (others => 'X'); -- umft_gpio_bus_signal
			umft_wr_n_pin                   : out   std_logic;                                         -- umft_wr_n_signal
			umft_rd_n_pin                   : out   std_logic;                                         -- umft_rd_n_signal
			umft_oe_n_pin                   : out   std_logic;                                         -- umft_oe_n_signal
			umft_siwu_n_pin                 : out   std_logic;                                         -- umft_siwu_n_signal
			avalon_slave_config_address     : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- address
			avalon_slave_config_write       : in    std_logic                      := 'X';             -- write
			avalon_slave_config_read        : in    std_logic                      := 'X';             -- read
			avalon_slave_config_readdata    : out   std_logic_vector(31 downto 0);                     -- readdata
			avalon_slave_config_writedata   : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			avalon_slave_config_waitrequest : out   std_logic;                                         -- waitrequest
			avalon_slave_config_byteenable  : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			avalon_slave_data_address       : in    std_logic_vector(20 downto 0)  := (others => 'X'); -- address
			avalon_slave_data_write         : in    std_logic                      := 'X';             -- write
			avalon_slave_data_read          : in    std_logic                      := 'X';             -- read
			avalon_slave_data_writedata     : in    std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			avalon_slave_data_readdata      : out   std_logic_vector(255 downto 0);                    -- readdata
			avalon_slave_data_waitrequest   : out   std_logic;                                         -- waitrequest
			ftdi_interrupt_sender_irq       : out   std_logic                                          -- irq
		);
	end component ftdi_usb3_top;

	component SEVEN_SEG_TOP is
		port (
			AVALON_SLAVE_ADDRESS   : in  std_logic                     := 'X';             -- address
			AVALON_SLAVE_WRITEDATA : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			AVALON_SLAVE_WRITE     : in  std_logic                     := 'X';             -- write
			CLK                    : in  std_logic                     := 'X';             -- clk
			RST                    : in  std_logic                     := 'X';             -- reset
			SEVEN_SEG_DSP0_OUT     : out std_logic_vector(7 downto 0);                     -- ssdp0
			SEVEN_SEG_DSP1_OUT     : out std_logic_vector(7 downto 0)                      -- ssdp1
		);
	end component SEVEN_SEG_TOP;

	component MebX_Qsys_Project_csense_adc_fo is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component MebX_Qsys_Project_csense_adc_fo;

	component MebX_Qsys_Project_csense_cs_n is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(1 downto 0)                      -- export
		);
	end component MebX_Qsys_Project_csense_cs_n;

	component MebX_Qsys_Project_csense_sdo is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component MebX_Qsys_Project_csense_sdo;

	component altera_address_span_extender is
		generic (
			DATA_WIDTH           : integer                       := 32;
			BYTEENABLE_WIDTH     : integer                       := 4;
			MASTER_ADDRESS_WIDTH : integer                       := 32;
			SLAVE_ADDRESS_WIDTH  : integer                       := 16;
			SLAVE_ADDRESS_SHIFT  : integer                       := 2;
			BURSTCOUNT_WIDTH     : integer                       := 1;
			CNTL_ADDRESS_WIDTH   : integer                       := 1;
			SUB_WINDOW_COUNT     : integer                       := 1;
			MASTER_ADDRESS_DEF   : std_logic_vector(63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000"
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			avs_s0_address       : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			avs_s0_read          : in  std_logic                     := 'X';             -- read
			avs_s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avs_s0_write         : in  std_logic                     := 'X';             -- write
			avs_s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_s0_readdatavalid : out std_logic;                                        -- readdatavalid
			avs_s0_waitrequest   : out std_logic;                                        -- waitrequest
			avs_s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_s0_burstcount    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			avm_m0_address       : out std_logic_vector(31 downto 0);                    -- address
			avm_m0_read          : out std_logic;                                        -- read
			avm_m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			avm_m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_m0_write         : out std_logic;                                        -- write
			avm_m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			avm_m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			avm_m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			avm_m0_burstcount    : out std_logic_vector(7 downto 0);                     -- burstcount
			avs_cntl_read        : in  std_logic                     := 'X';             -- read
			avs_cntl_readdata    : out std_logic_vector(63 downto 0);                    -- readdata
			avs_cntl_write       : in  std_logic                     := 'X';             -- write
			avs_cntl_writedata   : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			avs_cntl_byteenable  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			avs_cntl_address     : in  std_logic_vector(0 downto 0)  := (others => 'X')  -- address
		);
	end component altera_address_span_extender;

	component MebX_Qsys_Project_dma_comm_1_left is
		port (
			mm_read_address              : out std_logic_vector(31 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_read_readdata             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_write_address             : out std_logic_vector(32 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_write_writedata           : out std_logic_vector(255 downto 0);                    -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic                                          -- irq
		);
	end component MebX_Qsys_Project_dma_comm_1_left;

	component MebX_Qsys_Project_dma_comm_1_right is
		port (
			mm_read_address              : out std_logic_vector(31 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_read_readdata             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_write_address             : out std_logic_vector(32 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_write_writedata           : out std_logic_vector(255 downto 0);                    -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic                                          -- irq
		);
	end component MebX_Qsys_Project_dma_comm_1_right;

	component MebX_Qsys_Project_dma_comm_2_left is
		port (
			mm_read_address              : out std_logic_vector(31 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_read_readdata             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_write_address             : out std_logic_vector(32 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_write_writedata           : out std_logic_vector(255 downto 0);                    -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic                                          -- irq
		);
	end component MebX_Qsys_Project_dma_comm_2_left;

	component MebX_Qsys_Project_dma_comm_2_right is
		port (
			mm_read_address              : out std_logic_vector(31 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_read_readdata             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_write_address             : out std_logic_vector(32 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_write_writedata           : out std_logic_vector(255 downto 0);                    -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic                                          -- irq
		);
	end component MebX_Qsys_Project_dma_comm_2_right;

	component MebX_Qsys_Project_dma_comm_3_left is
		port (
			mm_read_address              : out std_logic_vector(31 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_read_readdata             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_write_address             : out std_logic_vector(32 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_write_writedata           : out std_logic_vector(255 downto 0);                    -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic                                          -- irq
		);
	end component MebX_Qsys_Project_dma_comm_3_left;

	component MebX_Qsys_Project_dma_comm_3_right is
		port (
			mm_read_address              : out std_logic_vector(31 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_read_readdata             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_write_address             : out std_logic_vector(32 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_write_writedata           : out std_logic_vector(255 downto 0);                    -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic                                          -- irq
		);
	end component MebX_Qsys_Project_dma_comm_3_right;

	component MebX_Qsys_Project_dma_comm_4_left is
		port (
			mm_read_address              : out std_logic_vector(31 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_read_readdata             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_write_address             : out std_logic_vector(32 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_write_writedata           : out std_logic_vector(255 downto 0);                    -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic                                          -- irq
		);
	end component MebX_Qsys_Project_dma_comm_4_left;

	component MebX_Qsys_Project_dma_comm_4_right is
		port (
			mm_read_address              : out std_logic_vector(31 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_read_readdata             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_write_address             : out std_logic_vector(32 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_write_writedata           : out std_logic_vector(255 downto 0);                    -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic                                          -- irq
		);
	end component MebX_Qsys_Project_dma_comm_4_right;

	component MebX_Qsys_Project_dma_comm_5_left is
		port (
			mm_read_address              : out std_logic_vector(31 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_read_readdata             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_write_address             : out std_logic_vector(32 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_write_writedata           : out std_logic_vector(255 downto 0);                    -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic                                          -- irq
		);
	end component MebX_Qsys_Project_dma_comm_5_left;

	component MebX_Qsys_Project_dma_comm_5_right is
		port (
			mm_read_address              : out std_logic_vector(31 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_read_readdata             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_write_address             : out std_logic_vector(32 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_write_writedata           : out std_logic_vector(255 downto 0);                    -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic                                          -- irq
		);
	end component MebX_Qsys_Project_dma_comm_5_right;

	component MebX_Qsys_Project_dma_comm_6_left is
		port (
			mm_read_address              : out std_logic_vector(31 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_read_readdata             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_write_address             : out std_logic_vector(32 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_write_writedata           : out std_logic_vector(255 downto 0);                    -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic                                          -- irq
		);
	end component MebX_Qsys_Project_dma_comm_6_left;

	component MebX_Qsys_Project_dma_comm_6_right is
		port (
			mm_read_address              : out std_logic_vector(31 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_read_readdata             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_write_address             : out std_logic_vector(32 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_write_writedata           : out std_logic_vector(255 downto 0);                    -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic                                          -- irq
		);
	end component MebX_Qsys_Project_dma_comm_6_right;

	component MebX_Qsys_Project_dma_ftdi_usb3 is
		port (
			mm_read_address              : out std_logic_vector(33 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_read_readdata             : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_write_address             : out std_logic_vector(31 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(31 downto 0);                     -- byteenable
			mm_write_writedata           : out std_logic_vector(255 downto 0);                    -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic                                          -- irq
		);
	end component MebX_Qsys_Project_dma_ftdi_usb3;

	component MebX_Qsys_Project_ext_flash is
		generic (
			TCM_ADDRESS_W                  : integer := 30;
			TCM_DATA_W                     : integer := 32;
			TCM_BYTEENABLE_W               : integer := 4;
			TCM_READ_WAIT                  : integer := 1;
			TCM_WRITE_WAIT                 : integer := 0;
			TCM_SETUP_WAIT                 : integer := 0;
			TCM_DATA_HOLD                  : integer := 0;
			TCM_TURNAROUND_TIME            : integer := 2;
			TCM_TIMING_UNITS               : integer := 1;
			TCM_READLATENCY                : integer := 2;
			TCM_SYMBOLS_PER_WORD           : integer := 4;
			USE_READDATA                   : integer := 1;
			USE_WRITEDATA                  : integer := 1;
			USE_READ                       : integer := 1;
			USE_WRITE                      : integer := 1;
			USE_BYTEENABLE                 : integer := 1;
			USE_CHIPSELECT                 : integer := 0;
			USE_LOCK                       : integer := 0;
			USE_ADDRESS                    : integer := 1;
			USE_WAITREQUEST                : integer := 0;
			USE_WRITEBYTEENABLE            : integer := 0;
			USE_OUTPUTENABLE               : integer := 0;
			USE_RESETREQUEST               : integer := 0;
			USE_IRQ                        : integer := 0;
			USE_RESET_OUTPUT               : integer := 0;
			ACTIVE_LOW_READ                : integer := 0;
			ACTIVE_LOW_LOCK                : integer := 0;
			ACTIVE_LOW_WRITE               : integer := 0;
			ACTIVE_LOW_CHIPSELECT          : integer := 0;
			ACTIVE_LOW_BYTEENABLE          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE        : integer := 0;
			ACTIVE_LOW_WRITEBYTEENABLE     : integer := 0;
			ACTIVE_LOW_WAITREQUEST         : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER       : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			reset_reset          : in  std_logic                     := 'X';             -- reset
			uas_address          : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			uas_burstcount       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uas_read             : in  std_logic                     := 'X';             -- read
			uas_write            : in  std_logic                     := 'X';             -- write
			uas_waitrequest      : out std_logic;                                        -- waitrequest
			uas_readdatavalid    : out std_logic;                                        -- readdatavalid
			uas_byteenable       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uas_readdata         : out std_logic_vector(15 downto 0);                    -- readdata
			uas_writedata        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uas_lock             : in  std_logic                     := 'X';             -- lock
			uas_debugaccess      : in  std_logic                     := 'X';             -- debugaccess
			tcm_write_n_out      : out std_logic;                                        -- write_n_out
			tcm_read_n_out       : out std_logic;                                        -- read_n_out
			tcm_chipselect_n_out : out std_logic;                                        -- chipselect_n_out
			tcm_request          : out std_logic;                                        -- request
			tcm_grant            : in  std_logic                     := 'X';             -- grant
			tcm_address_out      : out std_logic_vector(25 downto 0);                    -- address_out
			tcm_data_out         : out std_logic_vector(15 downto 0);                    -- data_out
			tcm_data_outen       : out std_logic;                                        -- data_outen
			tcm_data_in          : in  std_logic_vector(15 downto 0) := (others => 'X')  -- data_in
		);
	end component MebX_Qsys_Project_ext_flash;

	component MebX_Qsys_Project_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component MebX_Qsys_Project_jtag_uart_0;

	component MebX_Qsys_Project_m1_ddr2_i2c_sda is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic                     := 'X'              -- export
		);
	end component MebX_Qsys_Project_m1_ddr2_i2c_sda;

	component MebX_Qsys_Project_m1_ddr2_memory is
		port (
			pll_ref_clk        : in    std_logic                      := 'X';             -- clk
			global_reset_n     : in    std_logic                      := 'X';             -- reset_n
			soft_reset_n       : in    std_logic                      := 'X';             -- reset_n
			afi_clk            : out   std_logic;                                         -- clk
			afi_half_clk       : out   std_logic;                                         -- clk
			afi_reset_n        : out   std_logic;                                         -- reset_n
			afi_reset_export_n : out   std_logic;                                         -- reset_n
			mem_a              : out   std_logic_vector(13 downto 0);                     -- mem_a
			mem_ba             : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck             : out   std_logic_vector(1 downto 0);                      -- mem_ck
			mem_ck_n           : out   std_logic_vector(1 downto 0);                      -- mem_ck_n
			mem_cke            : out   std_logic_vector(1 downto 0);                      -- mem_cke
			mem_cs_n           : out   std_logic_vector(1 downto 0);                      -- mem_cs_n
			mem_dm             : out   std_logic_vector(7 downto 0);                      -- mem_dm
			mem_ras_n          : out   std_logic_vector(0 downto 0);                      -- mem_ras_n
			mem_cas_n          : out   std_logic_vector(0 downto 0);                      -- mem_cas_n
			mem_we_n           : out   std_logic_vector(0 downto 0);                      -- mem_we_n
			mem_dq             : inout std_logic_vector(63 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs            : inout std_logic_vector(7 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n          : inout std_logic_vector(7 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt            : out   std_logic_vector(1 downto 0);                      -- mem_odt
			avl_ready          : out   std_logic;                                         -- waitrequest_n
			avl_burstbegin     : in    std_logic                      := 'X';             -- beginbursttransfer
			avl_addr           : in    std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			avl_rdata_valid    : out   std_logic;                                         -- readdatavalid
			avl_rdata          : out   std_logic_vector(255 downto 0);                    -- readdata
			avl_wdata          : in    std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			avl_be             : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req       : in    std_logic                      := 'X';             -- read
			avl_write_req      : in    std_logic                      := 'X';             -- write
			avl_size           : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- burstcount
			local_init_done    : out   std_logic;                                         -- local_init_done
			local_cal_success  : out   std_logic;                                         -- local_cal_success
			local_cal_fail     : out   std_logic;                                         -- local_cal_fail
			oct_rdn            : in    std_logic                      := 'X';             -- rdn
			oct_rup            : in    std_logic                      := 'X'              -- rup
		);
	end component MebX_Qsys_Project_m1_ddr2_memory;

	component MebX_Qsys_Project_m2_ddr2_memory is
		port (
			pll_ref_clk               : in    std_logic                      := 'X';             -- clk
			global_reset_n            : in    std_logic                      := 'X';             -- reset_n
			soft_reset_n              : in    std_logic                      := 'X';             -- reset_n
			afi_clk                   : out   std_logic;                                         -- clk
			afi_half_clk              : out   std_logic;                                         -- clk
			afi_reset_n               : out   std_logic;                                         -- reset_n
			afi_reset_export_n        : out   std_logic;                                         -- reset_n
			mem_a                     : out   std_logic_vector(13 downto 0);                     -- mem_a
			mem_ba                    : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck                    : out   std_logic_vector(1 downto 0);                      -- mem_ck
			mem_ck_n                  : out   std_logic_vector(1 downto 0);                      -- mem_ck_n
			mem_cke                   : out   std_logic_vector(1 downto 0);                      -- mem_cke
			mem_cs_n                  : out   std_logic_vector(1 downto 0);                      -- mem_cs_n
			mem_dm                    : out   std_logic_vector(7 downto 0);                      -- mem_dm
			mem_ras_n                 : out   std_logic_vector(0 downto 0);                      -- mem_ras_n
			mem_cas_n                 : out   std_logic_vector(0 downto 0);                      -- mem_cas_n
			mem_we_n                  : out   std_logic_vector(0 downto 0);                      -- mem_we_n
			mem_dq                    : inout std_logic_vector(63 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs                   : inout std_logic_vector(7 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n                 : inout std_logic_vector(7 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt                   : out   std_logic_vector(1 downto 0);                      -- mem_odt
			avl_ready                 : out   std_logic;                                         -- waitrequest_n
			avl_burstbegin            : in    std_logic                      := 'X';             -- beginbursttransfer
			avl_addr                  : in    std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			avl_rdata_valid           : out   std_logic;                                         -- readdatavalid
			avl_rdata                 : out   std_logic_vector(255 downto 0);                    -- readdata
			avl_wdata                 : in    std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			avl_be                    : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req              : in    std_logic                      := 'X';             -- read
			avl_write_req             : in    std_logic                      := 'X';             -- write
			avl_size                  : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- burstcount
			local_init_done           : out   std_logic;                                         -- local_init_done
			local_cal_success         : out   std_logic;                                         -- local_cal_success
			local_cal_fail            : out   std_logic;                                         -- local_cal_fail
			oct_rdn                   : in    std_logic                      := 'X';             -- rdn
			oct_rup                   : in    std_logic                      := 'X';             -- rup
			pll_mem_clk               : out   std_logic;                                         -- pll_mem_clk
			pll_write_clk             : out   std_logic;                                         -- pll_write_clk
			pll_locked                : out   std_logic;                                         -- pll_locked
			pll_write_clk_pre_phy_clk : out   std_logic;                                         -- pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk          : out   std_logic;                                         -- pll_addr_cmd_clk
			pll_avl_clk               : out   std_logic;                                         -- pll_avl_clk
			pll_config_clk            : out   std_logic;                                         -- pll_config_clk
			dll_pll_locked            : in    std_logic                      := 'X';             -- dll_pll_locked
			dll_delayctrl             : out   std_logic_vector(5 downto 0)                       -- dll_delayctrl
		);
	end component MebX_Qsys_Project_m2_ddr2_memory;

	component MebX_Qsys_Project_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(31 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(31 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_burstcount                        : out std_logic_vector(3 downto 0);                     -- burstcount
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component MebX_Qsys_Project_nios2_gen2_0;

	component MebX_Qsys_Project_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component MebX_Qsys_Project_onchip_memory;

	component MebX_Qsys_Project_pio_BUTTON is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component MebX_Qsys_Project_pio_BUTTON;

	component MebX_Qsys_Project_pio_DIP is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component MebX_Qsys_Project_pio_DIP;

	component MebX_Qsys_Project_pio_EXT is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component MebX_Qsys_Project_pio_EXT;

	component MebX_Qsys_Project_pio_LED is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component MebX_Qsys_Project_pio_LED;

	component MebX_Qsys_Project_pio_LED_painel is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(20 downto 0)                     -- export
		);
	end component MebX_Qsys_Project_pio_LED_painel;

	component MebX_Qsys_Project_pio_ctrl_io_lvds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component MebX_Qsys_Project_pio_ctrl_io_lvds;

	component nrme_rmap_memory_nfee_area_top is
		port (
			reset_i                           : in  std_logic                     := 'X';             -- reset
			clk_100_i                         : in  std_logic                     := 'X';             -- clk
			avs_0_rmap_address_i              : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			avs_0_rmap_write_i                : in  std_logic                     := 'X';             -- write
			avs_0_rmap_read_i                 : in  std_logic                     := 'X';             -- read
			avs_0_rmap_readdata_o             : out std_logic_vector(31 downto 0);                    -- readdata
			avs_0_rmap_writedata_i            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_0_rmap_waitrequest_o          : out std_logic;                                        -- waitrequest
			avs_0_rmap_byteenable_i           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			fee_0_rmap_wr_address_i           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			fee_0_rmap_write_i                : in  std_logic                     := 'X';             -- write_signal
			fee_0_rmap_writedata_i            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			fee_0_rmap_rd_address_i           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			fee_0_rmap_read_i                 : in  std_logic                     := 'X';             -- read_signal
			fee_0_rmap_wr_waitrequest_o       : out std_logic;                                        -- wr_waitrequest_signal
			fee_0_rmap_readdata_o             : out std_logic_vector(7 downto 0);                     -- readdata_signal
			fee_0_rmap_rd_waitrequest_o       : out std_logic;                                        -- rd_waitrequest_signal
			fee_1_rmap_wr_address_i           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wr_address_signal
			fee_1_rmap_write_i                : in  std_logic                     := 'X';             -- write_signal
			fee_1_rmap_writedata_i            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata_signal
			fee_1_rmap_rd_address_i           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rd_address_signal
			fee_1_rmap_read_i                 : in  std_logic                     := 'X';             -- read_signal
			fee_1_rmap_wr_waitrequest_o       : out std_logic;                                        -- wr_waitrequest_signal
			fee_1_rmap_readdata_o             : out std_logic_vector(7 downto 0);                     -- readdata_signal
			fee_1_rmap_rd_waitrequest_o       : out std_logic;                                        -- rd_waitrequest_signal
			channel_hk_timecode_control_i     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- timecode_control_signal
			channel_hk_timecode_time_i        : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- timecode_time_signal
			channel_hk_rmap_target_status_i   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- rmap_target_status_signal
			channel_hk_rmap_target_indicate_i : in  std_logic                     := 'X';             -- rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_i  : in  std_logic                     := 'X';             -- spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_i  : in  std_logic                     := 'X';             -- spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_i  : in  std_logic                     := 'X';             -- spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_i  : in  std_logic                     := 'X';             -- spw_link_disconnect_signal
			channel_hk_spw_link_running_i     : in  std_logic                     := 'X';             -- spw_link_running_signal
			channel_hk_frame_counter_i        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- frame_counter_signal
			channel_hk_frame_number_i         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- frame_number_signal
			avm_rmap_readdata_i               : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			avm_rmap_waitrequest_i            : in  std_logic                     := 'X';             -- waitrequest
			avm_rmap_address_o                : out std_logic_vector(63 downto 0);                    -- address
			avm_rmap_read_o                   : out std_logic;                                        -- read
			avm_rmap_write_o                  : out std_logic;                                        -- write
			avm_rmap_writedata_o              : out std_logic_vector(7 downto 0);                     -- writedata
			channel_win_mem_addr_offset_i     : in  std_logic_vector(63 downto 0) := (others => 'X')  -- win_mem_addr_offset_signal
		);
	end component nrme_rmap_memory_nfee_area_top;

	component MebX_Qsys_Project_rs232_uart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component MebX_Qsys_Project_rs232_uart;

	component rst_controller_top is
		port (
			clock_sink_clk                          : in  std_logic                     := 'X';             -- clk
			reset_sink_reset                        : in  std_logic                     := 'X';             -- reset
			reset_source_ftdi_reset                 : out std_logic;                                        -- reset
			reset_source_sync_reset                 : out std_logic;                                        -- reset
			reset_source_rs232_reset                : out std_logic;                                        -- reset
			reset_source_sd_card_reset              : out std_logic;                                        -- reset
			reset_source_comm_ch8_reset             : out std_logic;                                        -- reset
			reset_source_comm_ch7_reset             : out std_logic;                                        -- reset
			reset_source_comm_ch6_reset             : out std_logic;                                        -- reset
			reset_source_comm_ch5_reset             : out std_logic;                                        -- reset
			reset_source_comm_ch4_reset             : out std_logic;                                        -- reset
			reset_source_comm_ch3_reset             : out std_logic;                                        -- reset
			reset_source_comm_ch2_reset             : out std_logic;                                        -- reset
			reset_source_comm_ch1_reset             : out std_logic;                                        -- reset
			avalon_slave_rst_controller_address     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			avalon_slave_rst_controller_write       : in  std_logic                     := 'X';             -- write
			avalon_slave_rst_controller_read        : in  std_logic                     := 'X';             -- read
			avalon_slave_rst_controller_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalon_slave_rst_controller_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avalon_slave_rst_controller_waitrequest : out std_logic;                                        -- waitrequest
			simucam_reset_signal                    : out std_logic;                                        -- t_simucam_reset_signal
			reset_input_signal                      : in  std_logic                     := 'X'              -- t_reset_input_signal
		);
	end component rst_controller_top;

	component sync_ent is
		generic (
			g_SYNC_IRQ_NUMBER     : natural := 0;
			g_PRE_SYNC_IRQ_NUMBER : natural := 0
		);
		port (
			clock_sink_clk_i                : in  std_logic                     := 'X';             -- clk
			reset_sink_reset_i              : in  std_logic                     := 'X';             -- reset
			avalon_slave_address_i          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			avalon_slave_read_i             : in  std_logic                     := 'X';             -- read
			avalon_slave_write_i            : in  std_logic                     := 'X';             -- write
			avalon_slave_writedata_i        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalon_slave_byteenable_i       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avalon_slave_readdata_o         : out std_logic_vector(31 downto 0);                    -- readdata
			avalon_slave_waitrequest_o      : out std_logic;                                        -- waitrequest
			conduit_sync_signal_syncin_i    : in  std_logic                     := 'X';             -- conduit
			conduit_sync_signal_spw1_o      : out std_logic;                                        -- conduit
			conduit_sync_signal_spw2_o      : out std_logic;                                        -- conduit
			conduit_sync_signal_spw3_o      : out std_logic;                                        -- conduit
			conduit_sync_signal_spw4_o      : out std_logic;                                        -- conduit
			conduit_sync_signal_spw5_o      : out std_logic;                                        -- conduit
			conduit_sync_signal_spw6_o      : out std_logic;                                        -- conduit
			conduit_sync_signal_spw7_o      : out std_logic;                                        -- conduit
			conduit_sync_signal_spw8_o      : out std_logic;                                        -- conduit
			conduit_sync_signal_syncout_o   : out std_logic;                                        -- conduit
			sync_interrupt_sender_irq_o     : out std_logic;                                        -- irq
			pre_sync_interrupt_sender_irq_o : out std_logic                                         -- irq
		);
	end component sync_ent;

	component MebX_Qsys_Project_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component MebX_Qsys_Project_sysid_qsys;

	component MebX_Qsys_Project_timer_1ms is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			timeout_pulse : out std_logic                                         -- export
		);
	end component MebX_Qsys_Project_timer_1ms;

	component MebX_Qsys_Project_timer_1us is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			timeout_pulse : out std_logic                                         -- export
		);
	end component MebX_Qsys_Project_timer_1us;

	component MebX_Qsys_Project_tristate_conduit_bridge_0 is
		port (
			clk                      : in    std_logic                     := 'X';             -- clk
			reset                    : in    std_logic                     := 'X';             -- reset
			request                  : in    std_logic                     := 'X';             -- request
			grant                    : out   std_logic;                                        -- grant
			tcs_tcm_address_out      : in    std_logic_vector(25 downto 0) := (others => 'X'); -- address_out
			tcs_tcm_read_n_out       : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- read_n_out
			tcs_tcm_write_n_out      : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_out
			tcs_tcm_data_out         : in    std_logic_vector(15 downto 0) := (others => 'X'); -- data_out
			tcs_tcm_data_outen       : in    std_logic                     := 'X';             -- data_outen
			tcs_tcm_data_in          : out   std_logic_vector(15 downto 0);                    -- data_in
			tcs_tcm_chipselect_n_out : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- chipselect_n_out
			tcm_address_out          : out   std_logic_vector(25 downto 0);                    -- tcm_address_out
			tcm_read_n_out           : out   std_logic_vector(0 downto 0);                     -- tcm_read_n_out
			tcm_write_n_out          : out   std_logic_vector(0 downto 0);                     -- tcm_write_n_out
			tcm_data_out             : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			tcm_chipselect_n_out     : out   std_logic_vector(0 downto 0)                      -- tcm_chipselect_n_out
		);
	end component MebX_Qsys_Project_tristate_conduit_bridge_0;

	component MebX_Qsys_Project_mm_interconnect_0 is
		port (
			clk_100_clk_clk                                                 : in  std_logic                      := 'X';             -- clk
			m2_ddr2_memory_afi_clk_clk                                      : in  std_logic                      := 'X';             -- clk
			m2_ddr2_memory_afi_half_clk_clk                                 : in  std_logic                      := 'X';             -- clk
			ddr2_address_span_extender_reset_reset_bridge_in_reset_reset    : in  std_logic                      := 'X';             -- reset
			m1_clock_bridge_s0_reset_reset_bridge_in_reset_reset            : in  std_logic                      := 'X';             -- reset
			m2_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			m2_ddr2_memory_soft_reset_reset_bridge_in_reset_reset           : in  std_logic                      := 'X';             -- reset
			rmap_mem_nfee_comm_1_reset_sink_reset_bridge_in_reset_reset     : in  std_logic                      := 'X';             -- reset
			rmap_mem_nfee_comm_2_reset_sink_reset_bridge_in_reset_reset     : in  std_logic                      := 'X';             -- reset
			rmap_mem_nfee_comm_3_reset_sink_reset_bridge_in_reset_reset     : in  std_logic                      := 'X';             -- reset
			rmap_mem_nfee_comm_4_reset_sink_reset_bridge_in_reset_reset     : in  std_logic                      := 'X';             -- reset
			rmap_mem_nfee_comm_5_reset_sink_reset_bridge_in_reset_reset     : in  std_logic                      := 'X';             -- reset
			rmap_mem_nfee_comm_6_reset_sink_reset_bridge_in_reset_reset     : in  std_logic                      := 'X';             -- reset
			ddr2_address_span_extender_expanded_master_address              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			ddr2_address_span_extender_expanded_master_waitrequest          : out std_logic;                                         -- waitrequest
			ddr2_address_span_extender_expanded_master_burstcount           : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- burstcount
			ddr2_address_span_extender_expanded_master_byteenable           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			ddr2_address_span_extender_expanded_master_read                 : in  std_logic                      := 'X';             -- read
			ddr2_address_span_extender_expanded_master_readdata             : out std_logic_vector(31 downto 0);                     -- readdata
			ddr2_address_span_extender_expanded_master_readdatavalid        : out std_logic;                                         -- readdatavalid
			ddr2_address_span_extender_expanded_master_write                : in  std_logic                      := 'X';             -- write
			ddr2_address_span_extender_expanded_master_writedata            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			dma_comm_1_left_mm_read_address                                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			dma_comm_1_left_mm_read_waitrequest                             : out std_logic;                                         -- waitrequest
			dma_comm_1_left_mm_read_byteenable                              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_1_left_mm_read_read                                    : in  std_logic                      := 'X';             -- read
			dma_comm_1_left_mm_read_readdata                                : out std_logic_vector(255 downto 0);                    -- readdata
			dma_comm_1_left_mm_read_readdatavalid                           : out std_logic;                                         -- readdatavalid
			dma_comm_1_right_mm_read_address                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			dma_comm_1_right_mm_read_waitrequest                            : out std_logic;                                         -- waitrequest
			dma_comm_1_right_mm_read_byteenable                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_1_right_mm_read_read                                   : in  std_logic                      := 'X';             -- read
			dma_comm_1_right_mm_read_readdata                               : out std_logic_vector(255 downto 0);                    -- readdata
			dma_comm_1_right_mm_read_readdatavalid                          : out std_logic;                                         -- readdatavalid
			dma_comm_2_left_mm_read_address                                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			dma_comm_2_left_mm_read_waitrequest                             : out std_logic;                                         -- waitrequest
			dma_comm_2_left_mm_read_byteenable                              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_2_left_mm_read_read                                    : in  std_logic                      := 'X';             -- read
			dma_comm_2_left_mm_read_readdata                                : out std_logic_vector(255 downto 0);                    -- readdata
			dma_comm_2_left_mm_read_readdatavalid                           : out std_logic;                                         -- readdatavalid
			dma_comm_2_right_mm_read_address                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			dma_comm_2_right_mm_read_waitrequest                            : out std_logic;                                         -- waitrequest
			dma_comm_2_right_mm_read_byteenable                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_2_right_mm_read_read                                   : in  std_logic                      := 'X';             -- read
			dma_comm_2_right_mm_read_readdata                               : out std_logic_vector(255 downto 0);                    -- readdata
			dma_comm_2_right_mm_read_readdatavalid                          : out std_logic;                                         -- readdatavalid
			dma_comm_3_left_mm_read_address                                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			dma_comm_3_left_mm_read_waitrequest                             : out std_logic;                                         -- waitrequest
			dma_comm_3_left_mm_read_byteenable                              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_3_left_mm_read_read                                    : in  std_logic                      := 'X';             -- read
			dma_comm_3_left_mm_read_readdata                                : out std_logic_vector(255 downto 0);                    -- readdata
			dma_comm_3_left_mm_read_readdatavalid                           : out std_logic;                                         -- readdatavalid
			dma_comm_3_right_mm_read_address                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			dma_comm_3_right_mm_read_waitrequest                            : out std_logic;                                         -- waitrequest
			dma_comm_3_right_mm_read_byteenable                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_3_right_mm_read_read                                   : in  std_logic                      := 'X';             -- read
			dma_comm_3_right_mm_read_readdata                               : out std_logic_vector(255 downto 0);                    -- readdata
			dma_comm_3_right_mm_read_readdatavalid                          : out std_logic;                                         -- readdatavalid
			dma_comm_4_left_mm_read_address                                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			dma_comm_4_left_mm_read_waitrequest                             : out std_logic;                                         -- waitrequest
			dma_comm_4_left_mm_read_byteenable                              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_4_left_mm_read_read                                    : in  std_logic                      := 'X';             -- read
			dma_comm_4_left_mm_read_readdata                                : out std_logic_vector(255 downto 0);                    -- readdata
			dma_comm_4_left_mm_read_readdatavalid                           : out std_logic;                                         -- readdatavalid
			dma_comm_4_right_mm_read_address                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			dma_comm_4_right_mm_read_waitrequest                            : out std_logic;                                         -- waitrequest
			dma_comm_4_right_mm_read_byteenable                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_4_right_mm_read_read                                   : in  std_logic                      := 'X';             -- read
			dma_comm_4_right_mm_read_readdata                               : out std_logic_vector(255 downto 0);                    -- readdata
			dma_comm_4_right_mm_read_readdatavalid                          : out std_logic;                                         -- readdatavalid
			dma_comm_5_left_mm_read_address                                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			dma_comm_5_left_mm_read_waitrequest                             : out std_logic;                                         -- waitrequest
			dma_comm_5_left_mm_read_byteenable                              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_5_left_mm_read_read                                    : in  std_logic                      := 'X';             -- read
			dma_comm_5_left_mm_read_readdata                                : out std_logic_vector(255 downto 0);                    -- readdata
			dma_comm_5_left_mm_read_readdatavalid                           : out std_logic;                                         -- readdatavalid
			dma_comm_5_right_mm_read_address                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			dma_comm_5_right_mm_read_waitrequest                            : out std_logic;                                         -- waitrequest
			dma_comm_5_right_mm_read_byteenable                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_5_right_mm_read_read                                   : in  std_logic                      := 'X';             -- read
			dma_comm_5_right_mm_read_readdata                               : out std_logic_vector(255 downto 0);                    -- readdata
			dma_comm_5_right_mm_read_readdatavalid                          : out std_logic;                                         -- readdatavalid
			dma_comm_6_left_mm_read_address                                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			dma_comm_6_left_mm_read_waitrequest                             : out std_logic;                                         -- waitrequest
			dma_comm_6_left_mm_read_byteenable                              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_6_left_mm_read_read                                    : in  std_logic                      := 'X';             -- read
			dma_comm_6_left_mm_read_readdata                                : out std_logic_vector(255 downto 0);                    -- readdata
			dma_comm_6_left_mm_read_readdatavalid                           : out std_logic;                                         -- readdatavalid
			dma_comm_6_right_mm_read_address                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			dma_comm_6_right_mm_read_waitrequest                            : out std_logic;                                         -- waitrequest
			dma_comm_6_right_mm_read_byteenable                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_6_right_mm_read_read                                   : in  std_logic                      := 'X';             -- read
			dma_comm_6_right_mm_read_readdata                               : out std_logic_vector(255 downto 0);                    -- readdata
			dma_comm_6_right_mm_read_readdatavalid                          : out std_logic;                                         -- readdatavalid
			dma_ftdi_usb3_mm_write_address                                  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			dma_ftdi_usb3_mm_write_waitrequest                              : out std_logic;                                         -- waitrequest
			dma_ftdi_usb3_mm_write_byteenable                               : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_ftdi_usb3_mm_write_write                                    : in  std_logic                      := 'X';             -- write
			dma_ftdi_usb3_mm_write_writedata                                : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			rmap_mem_nfee_comm_1_avalon_mm_rmap_master_address              : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			rmap_mem_nfee_comm_1_avalon_mm_rmap_master_waitrequest          : out std_logic;                                         -- waitrequest
			rmap_mem_nfee_comm_1_avalon_mm_rmap_master_read                 : in  std_logic                      := 'X';             -- read
			rmap_mem_nfee_comm_1_avalon_mm_rmap_master_readdata             : out std_logic_vector(7 downto 0);                      -- readdata
			rmap_mem_nfee_comm_1_avalon_mm_rmap_master_write                : in  std_logic                      := 'X';             -- write
			rmap_mem_nfee_comm_1_avalon_mm_rmap_master_writedata            : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- writedata
			rmap_mem_nfee_comm_2_avalon_mm_rmap_master_address              : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			rmap_mem_nfee_comm_2_avalon_mm_rmap_master_waitrequest          : out std_logic;                                         -- waitrequest
			rmap_mem_nfee_comm_2_avalon_mm_rmap_master_read                 : in  std_logic                      := 'X';             -- read
			rmap_mem_nfee_comm_2_avalon_mm_rmap_master_readdata             : out std_logic_vector(7 downto 0);                      -- readdata
			rmap_mem_nfee_comm_2_avalon_mm_rmap_master_write                : in  std_logic                      := 'X';             -- write
			rmap_mem_nfee_comm_2_avalon_mm_rmap_master_writedata            : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- writedata
			rmap_mem_nfee_comm_3_avalon_mm_rmap_master_address              : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			rmap_mem_nfee_comm_3_avalon_mm_rmap_master_waitrequest          : out std_logic;                                         -- waitrequest
			rmap_mem_nfee_comm_3_avalon_mm_rmap_master_read                 : in  std_logic                      := 'X';             -- read
			rmap_mem_nfee_comm_3_avalon_mm_rmap_master_readdata             : out std_logic_vector(7 downto 0);                      -- readdata
			rmap_mem_nfee_comm_3_avalon_mm_rmap_master_write                : in  std_logic                      := 'X';             -- write
			rmap_mem_nfee_comm_3_avalon_mm_rmap_master_writedata            : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- writedata
			rmap_mem_nfee_comm_4_avalon_mm_rmap_master_address              : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			rmap_mem_nfee_comm_4_avalon_mm_rmap_master_waitrequest          : out std_logic;                                         -- waitrequest
			rmap_mem_nfee_comm_4_avalon_mm_rmap_master_read                 : in  std_logic                      := 'X';             -- read
			rmap_mem_nfee_comm_4_avalon_mm_rmap_master_readdata             : out std_logic_vector(7 downto 0);                      -- readdata
			rmap_mem_nfee_comm_4_avalon_mm_rmap_master_write                : in  std_logic                      := 'X';             -- write
			rmap_mem_nfee_comm_4_avalon_mm_rmap_master_writedata            : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- writedata
			rmap_mem_nfee_comm_5_avalon_mm_rmap_master_address              : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			rmap_mem_nfee_comm_5_avalon_mm_rmap_master_waitrequest          : out std_logic;                                         -- waitrequest
			rmap_mem_nfee_comm_5_avalon_mm_rmap_master_read                 : in  std_logic                      := 'X';             -- read
			rmap_mem_nfee_comm_5_avalon_mm_rmap_master_readdata             : out std_logic_vector(7 downto 0);                      -- readdata
			rmap_mem_nfee_comm_5_avalon_mm_rmap_master_write                : in  std_logic                      := 'X';             -- write
			rmap_mem_nfee_comm_5_avalon_mm_rmap_master_writedata            : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- writedata
			rmap_mem_nfee_comm_6_avalon_mm_rmap_master_address              : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- address
			rmap_mem_nfee_comm_6_avalon_mm_rmap_master_waitrequest          : out std_logic;                                         -- waitrequest
			rmap_mem_nfee_comm_6_avalon_mm_rmap_master_read                 : in  std_logic                      := 'X';             -- read
			rmap_mem_nfee_comm_6_avalon_mm_rmap_master_readdata             : out std_logic_vector(7 downto 0);                      -- readdata
			rmap_mem_nfee_comm_6_avalon_mm_rmap_master_write                : in  std_logic                      := 'X';             -- write
			rmap_mem_nfee_comm_6_avalon_mm_rmap_master_writedata            : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- writedata
			m1_clock_bridge_s0_address                                      : out std_logic_vector(30 downto 0);                     -- address
			m1_clock_bridge_s0_write                                        : out std_logic;                                         -- write
			m1_clock_bridge_s0_read                                         : out std_logic;                                         -- read
			m1_clock_bridge_s0_readdata                                     : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			m1_clock_bridge_s0_writedata                                    : out std_logic_vector(255 downto 0);                    -- writedata
			m1_clock_bridge_s0_burstcount                                   : out std_logic_vector(2 downto 0);                      -- burstcount
			m1_clock_bridge_s0_byteenable                                   : out std_logic_vector(31 downto 0);                     -- byteenable
			m1_clock_bridge_s0_readdatavalid                                : in  std_logic                      := 'X';             -- readdatavalid
			m1_clock_bridge_s0_waitrequest                                  : in  std_logic                      := 'X';             -- waitrequest
			m1_clock_bridge_s0_debugaccess                                  : out std_logic;                                         -- debugaccess
			m2_ddr2_memory_avl_address                                      : out std_logic_vector(25 downto 0);                     -- address
			m2_ddr2_memory_avl_write                                        : out std_logic;                                         -- write
			m2_ddr2_memory_avl_read                                         : out std_logic;                                         -- read
			m2_ddr2_memory_avl_readdata                                     : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			m2_ddr2_memory_avl_writedata                                    : out std_logic_vector(255 downto 0);                    -- writedata
			m2_ddr2_memory_avl_beginbursttransfer                           : out std_logic;                                         -- beginbursttransfer
			m2_ddr2_memory_avl_burstcount                                   : out std_logic_vector(7 downto 0);                      -- burstcount
			m2_ddr2_memory_avl_byteenable                                   : out std_logic_vector(31 downto 0);                     -- byteenable
			m2_ddr2_memory_avl_readdatavalid                                : in  std_logic                      := 'X';             -- readdatavalid
			m2_ddr2_memory_avl_waitrequest                                  : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_0;

	component MebX_Qsys_Project_mm_interconnect_1 is
		port (
			clk_100_clk_clk                                             : in  std_logic                      := 'X';             -- clk
			ext_flash_reset_reset_bridge_in_reset_reset                 : in  std_logic                      := 'X';             -- reset
			jtag_uart_0_reset_reset_bridge_in_reset_reset               : in  std_logic                      := 'X';             -- reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset              : in  std_logic                      := 'X';             -- reset
			rmap_mem_nfee_comm_1_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			rmap_mem_nfee_comm_2_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			rmap_mem_nfee_comm_3_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			rmap_mem_nfee_comm_4_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			rmap_mem_nfee_comm_5_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			rmap_mem_nfee_comm_6_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			nios2_gen2_0_data_master_address                            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                        : out std_logic;                                         -- waitrequest
			nios2_gen2_0_data_master_byteenable                         : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                               : in  std_logic                      := 'X';             -- read
			nios2_gen2_0_data_master_readdata                           : out std_logic_vector(31 downto 0);                     -- readdata
			nios2_gen2_0_data_master_write                              : in  std_logic                      := 'X';             -- write
			nios2_gen2_0_data_master_writedata                          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                        : in  std_logic                      := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address                     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest                 : out std_logic;                                         -- waitrequest
			nios2_gen2_0_instruction_master_burstcount                  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			nios2_gen2_0_instruction_master_read                        : in  std_logic                      := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata                    : out std_logic_vector(31 downto 0);                     -- readdata
			nios2_gen2_0_instruction_master_readdatavalid               : out std_logic;                                         -- readdatavalid
			clock_bridge_afi_50_s0_address                              : out std_logic_vector(11 downto 0);                     -- address
			clock_bridge_afi_50_s0_write                                : out std_logic;                                         -- write
			clock_bridge_afi_50_s0_read                                 : out std_logic;                                         -- read
			clock_bridge_afi_50_s0_readdata                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			clock_bridge_afi_50_s0_writedata                            : out std_logic_vector(31 downto 0);                     -- writedata
			clock_bridge_afi_50_s0_burstcount                           : out std_logic_vector(0 downto 0);                      -- burstcount
			clock_bridge_afi_50_s0_byteenable                           : out std_logic_vector(3 downto 0);                      -- byteenable
			clock_bridge_afi_50_s0_readdatavalid                        : in  std_logic                      := 'X';             -- readdatavalid
			clock_bridge_afi_50_s0_waitrequest                          : in  std_logic                      := 'X';             -- waitrequest
			clock_bridge_afi_50_s0_debugaccess                          : out std_logic;                                         -- debugaccess
			COMM_Pedreiro_v1_01_A_avalon_slave_windowing_address        : out std_logic_vector(7 downto 0);                      -- address
			COMM_Pedreiro_v1_01_A_avalon_slave_windowing_write          : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_A_avalon_slave_windowing_read           : out std_logic;                                         -- read
			COMM_Pedreiro_v1_01_A_avalon_slave_windowing_readdata       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			COMM_Pedreiro_v1_01_A_avalon_slave_windowing_writedata      : out std_logic_vector(31 downto 0);                     -- writedata
			COMM_Pedreiro_v1_01_A_avalon_slave_windowing_byteenable     : out std_logic_vector(3 downto 0);                      -- byteenable
			COMM_Pedreiro_v1_01_A_avalon_slave_windowing_waitrequest    : in  std_logic                      := 'X';             -- waitrequest
			COMM_Pedreiro_v1_01_B_avalon_slave_windowing_address        : out std_logic_vector(7 downto 0);                      -- address
			COMM_Pedreiro_v1_01_B_avalon_slave_windowing_write          : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_B_avalon_slave_windowing_read           : out std_logic;                                         -- read
			COMM_Pedreiro_v1_01_B_avalon_slave_windowing_readdata       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			COMM_Pedreiro_v1_01_B_avalon_slave_windowing_writedata      : out std_logic_vector(31 downto 0);                     -- writedata
			COMM_Pedreiro_v1_01_B_avalon_slave_windowing_byteenable     : out std_logic_vector(3 downto 0);                      -- byteenable
			COMM_Pedreiro_v1_01_B_avalon_slave_windowing_waitrequest    : in  std_logic                      := 'X';             -- waitrequest
			COMM_Pedreiro_v1_01_C_avalon_slave_windowing_address        : out std_logic_vector(7 downto 0);                      -- address
			COMM_Pedreiro_v1_01_C_avalon_slave_windowing_write          : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_C_avalon_slave_windowing_read           : out std_logic;                                         -- read
			COMM_Pedreiro_v1_01_C_avalon_slave_windowing_readdata       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			COMM_Pedreiro_v1_01_C_avalon_slave_windowing_writedata      : out std_logic_vector(31 downto 0);                     -- writedata
			COMM_Pedreiro_v1_01_C_avalon_slave_windowing_byteenable     : out std_logic_vector(3 downto 0);                      -- byteenable
			COMM_Pedreiro_v1_01_C_avalon_slave_windowing_waitrequest    : in  std_logic                      := 'X';             -- waitrequest
			COMM_Pedreiro_v1_01_D_avalon_slave_windowing_address        : out std_logic_vector(7 downto 0);                      -- address
			COMM_Pedreiro_v1_01_D_avalon_slave_windowing_write          : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_D_avalon_slave_windowing_read           : out std_logic;                                         -- read
			COMM_Pedreiro_v1_01_D_avalon_slave_windowing_readdata       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			COMM_Pedreiro_v1_01_D_avalon_slave_windowing_writedata      : out std_logic_vector(31 downto 0);                     -- writedata
			COMM_Pedreiro_v1_01_D_avalon_slave_windowing_byteenable     : out std_logic_vector(3 downto 0);                      -- byteenable
			COMM_Pedreiro_v1_01_D_avalon_slave_windowing_waitrequest    : in  std_logic                      := 'X';             -- waitrequest
			COMM_Pedreiro_v1_01_E_avalon_slave_windowing_address        : out std_logic_vector(7 downto 0);                      -- address
			COMM_Pedreiro_v1_01_E_avalon_slave_windowing_write          : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_E_avalon_slave_windowing_read           : out std_logic;                                         -- read
			COMM_Pedreiro_v1_01_E_avalon_slave_windowing_readdata       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			COMM_Pedreiro_v1_01_E_avalon_slave_windowing_writedata      : out std_logic_vector(31 downto 0);                     -- writedata
			COMM_Pedreiro_v1_01_E_avalon_slave_windowing_byteenable     : out std_logic_vector(3 downto 0);                      -- byteenable
			COMM_Pedreiro_v1_01_E_avalon_slave_windowing_waitrequest    : in  std_logic                      := 'X';             -- waitrequest
			COMM_Pedreiro_v1_01_F_avalon_slave_windowing_address        : out std_logic_vector(7 downto 0);                      -- address
			COMM_Pedreiro_v1_01_F_avalon_slave_windowing_write          : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_F_avalon_slave_windowing_read           : out std_logic;                                         -- read
			COMM_Pedreiro_v1_01_F_avalon_slave_windowing_readdata       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			COMM_Pedreiro_v1_01_F_avalon_slave_windowing_writedata      : out std_logic_vector(31 downto 0);                     -- writedata
			COMM_Pedreiro_v1_01_F_avalon_slave_windowing_byteenable     : out std_logic_vector(3 downto 0);                      -- byteenable
			COMM_Pedreiro_v1_01_F_avalon_slave_windowing_waitrequest    : in  std_logic                      := 'X';             -- waitrequest
			ddr2_address_span_extender_cntl_write                       : out std_logic;                                         -- write
			ddr2_address_span_extender_cntl_read                        : out std_logic;                                         -- read
			ddr2_address_span_extender_cntl_readdata                    : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- readdata
			ddr2_address_span_extender_cntl_writedata                   : out std_logic_vector(63 downto 0);                     -- writedata
			ddr2_address_span_extender_cntl_byteenable                  : out std_logic_vector(7 downto 0);                      -- byteenable
			ddr2_address_span_extender_windowed_slave_address           : out std_logic_vector(28 downto 0);                     -- address
			ddr2_address_span_extender_windowed_slave_write             : out std_logic;                                         -- write
			ddr2_address_span_extender_windowed_slave_read              : out std_logic;                                         -- read
			ddr2_address_span_extender_windowed_slave_readdata          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			ddr2_address_span_extender_windowed_slave_writedata         : out std_logic_vector(31 downto 0);                     -- writedata
			ddr2_address_span_extender_windowed_slave_burstcount        : out std_logic_vector(7 downto 0);                      -- burstcount
			ddr2_address_span_extender_windowed_slave_byteenable        : out std_logic_vector(3 downto 0);                      -- byteenable
			ddr2_address_span_extender_windowed_slave_readdatavalid     : in  std_logic                      := 'X';             -- readdatavalid
			ddr2_address_span_extender_windowed_slave_waitrequest       : in  std_logic                      := 'X';             -- waitrequest
			dma_comm_1_left_csr_address                                 : out std_logic_vector(2 downto 0);                      -- address
			dma_comm_1_left_csr_write                                   : out std_logic;                                         -- write
			dma_comm_1_left_csr_read                                    : out std_logic;                                         -- read
			dma_comm_1_left_csr_readdata                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_comm_1_left_csr_writedata                               : out std_logic_vector(31 downto 0);                     -- writedata
			dma_comm_1_left_csr_byteenable                              : out std_logic_vector(3 downto 0);                      -- byteenable
			dma_comm_1_left_descriptor_slave_write                      : out std_logic;                                         -- write
			dma_comm_1_left_descriptor_slave_writedata                  : out std_logic_vector(255 downto 0);                    -- writedata
			dma_comm_1_left_descriptor_slave_byteenable                 : out std_logic_vector(31 downto 0);                     -- byteenable
			dma_comm_1_left_descriptor_slave_waitrequest                : in  std_logic                      := 'X';             -- waitrequest
			dma_comm_1_right_csr_address                                : out std_logic_vector(2 downto 0);                      -- address
			dma_comm_1_right_csr_write                                  : out std_logic;                                         -- write
			dma_comm_1_right_csr_read                                   : out std_logic;                                         -- read
			dma_comm_1_right_csr_readdata                               : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_comm_1_right_csr_writedata                              : out std_logic_vector(31 downto 0);                     -- writedata
			dma_comm_1_right_csr_byteenable                             : out std_logic_vector(3 downto 0);                      -- byteenable
			dma_comm_1_right_descriptor_slave_write                     : out std_logic;                                         -- write
			dma_comm_1_right_descriptor_slave_writedata                 : out std_logic_vector(255 downto 0);                    -- writedata
			dma_comm_1_right_descriptor_slave_byteenable                : out std_logic_vector(31 downto 0);                     -- byteenable
			dma_comm_1_right_descriptor_slave_waitrequest               : in  std_logic                      := 'X';             -- waitrequest
			dma_comm_2_left_csr_address                                 : out std_logic_vector(2 downto 0);                      -- address
			dma_comm_2_left_csr_write                                   : out std_logic;                                         -- write
			dma_comm_2_left_csr_read                                    : out std_logic;                                         -- read
			dma_comm_2_left_csr_readdata                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_comm_2_left_csr_writedata                               : out std_logic_vector(31 downto 0);                     -- writedata
			dma_comm_2_left_csr_byteenable                              : out std_logic_vector(3 downto 0);                      -- byteenable
			dma_comm_2_left_descriptor_slave_write                      : out std_logic;                                         -- write
			dma_comm_2_left_descriptor_slave_writedata                  : out std_logic_vector(255 downto 0);                    -- writedata
			dma_comm_2_left_descriptor_slave_byteenable                 : out std_logic_vector(31 downto 0);                     -- byteenable
			dma_comm_2_left_descriptor_slave_waitrequest                : in  std_logic                      := 'X';             -- waitrequest
			dma_comm_2_right_csr_address                                : out std_logic_vector(2 downto 0);                      -- address
			dma_comm_2_right_csr_write                                  : out std_logic;                                         -- write
			dma_comm_2_right_csr_read                                   : out std_logic;                                         -- read
			dma_comm_2_right_csr_readdata                               : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_comm_2_right_csr_writedata                              : out std_logic_vector(31 downto 0);                     -- writedata
			dma_comm_2_right_csr_byteenable                             : out std_logic_vector(3 downto 0);                      -- byteenable
			dma_comm_2_right_descriptor_slave_write                     : out std_logic;                                         -- write
			dma_comm_2_right_descriptor_slave_writedata                 : out std_logic_vector(255 downto 0);                    -- writedata
			dma_comm_2_right_descriptor_slave_byteenable                : out std_logic_vector(31 downto 0);                     -- byteenable
			dma_comm_2_right_descriptor_slave_waitrequest               : in  std_logic                      := 'X';             -- waitrequest
			dma_comm_3_left_csr_address                                 : out std_logic_vector(2 downto 0);                      -- address
			dma_comm_3_left_csr_write                                   : out std_logic;                                         -- write
			dma_comm_3_left_csr_read                                    : out std_logic;                                         -- read
			dma_comm_3_left_csr_readdata                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_comm_3_left_csr_writedata                               : out std_logic_vector(31 downto 0);                     -- writedata
			dma_comm_3_left_csr_byteenable                              : out std_logic_vector(3 downto 0);                      -- byteenable
			dma_comm_3_left_descriptor_slave_write                      : out std_logic;                                         -- write
			dma_comm_3_left_descriptor_slave_writedata                  : out std_logic_vector(255 downto 0);                    -- writedata
			dma_comm_3_left_descriptor_slave_byteenable                 : out std_logic_vector(31 downto 0);                     -- byteenable
			dma_comm_3_left_descriptor_slave_waitrequest                : in  std_logic                      := 'X';             -- waitrequest
			dma_comm_3_right_csr_address                                : out std_logic_vector(2 downto 0);                      -- address
			dma_comm_3_right_csr_write                                  : out std_logic;                                         -- write
			dma_comm_3_right_csr_read                                   : out std_logic;                                         -- read
			dma_comm_3_right_csr_readdata                               : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_comm_3_right_csr_writedata                              : out std_logic_vector(31 downto 0);                     -- writedata
			dma_comm_3_right_csr_byteenable                             : out std_logic_vector(3 downto 0);                      -- byteenable
			dma_comm_3_right_descriptor_slave_write                     : out std_logic;                                         -- write
			dma_comm_3_right_descriptor_slave_writedata                 : out std_logic_vector(255 downto 0);                    -- writedata
			dma_comm_3_right_descriptor_slave_byteenable                : out std_logic_vector(31 downto 0);                     -- byteenable
			dma_comm_3_right_descriptor_slave_waitrequest               : in  std_logic                      := 'X';             -- waitrequest
			dma_comm_4_left_csr_address                                 : out std_logic_vector(2 downto 0);                      -- address
			dma_comm_4_left_csr_write                                   : out std_logic;                                         -- write
			dma_comm_4_left_csr_read                                    : out std_logic;                                         -- read
			dma_comm_4_left_csr_readdata                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_comm_4_left_csr_writedata                               : out std_logic_vector(31 downto 0);                     -- writedata
			dma_comm_4_left_csr_byteenable                              : out std_logic_vector(3 downto 0);                      -- byteenable
			dma_comm_4_left_descriptor_slave_write                      : out std_logic;                                         -- write
			dma_comm_4_left_descriptor_slave_writedata                  : out std_logic_vector(255 downto 0);                    -- writedata
			dma_comm_4_left_descriptor_slave_byteenable                 : out std_logic_vector(31 downto 0);                     -- byteenable
			dma_comm_4_left_descriptor_slave_waitrequest                : in  std_logic                      := 'X';             -- waitrequest
			dma_comm_4_right_csr_address                                : out std_logic_vector(2 downto 0);                      -- address
			dma_comm_4_right_csr_write                                  : out std_logic;                                         -- write
			dma_comm_4_right_csr_read                                   : out std_logic;                                         -- read
			dma_comm_4_right_csr_readdata                               : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_comm_4_right_csr_writedata                              : out std_logic_vector(31 downto 0);                     -- writedata
			dma_comm_4_right_csr_byteenable                             : out std_logic_vector(3 downto 0);                      -- byteenable
			dma_comm_4_right_descriptor_slave_write                     : out std_logic;                                         -- write
			dma_comm_4_right_descriptor_slave_writedata                 : out std_logic_vector(255 downto 0);                    -- writedata
			dma_comm_4_right_descriptor_slave_byteenable                : out std_logic_vector(31 downto 0);                     -- byteenable
			dma_comm_4_right_descriptor_slave_waitrequest               : in  std_logic                      := 'X';             -- waitrequest
			dma_comm_5_left_csr_address                                 : out std_logic_vector(2 downto 0);                      -- address
			dma_comm_5_left_csr_write                                   : out std_logic;                                         -- write
			dma_comm_5_left_csr_read                                    : out std_logic;                                         -- read
			dma_comm_5_left_csr_readdata                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_comm_5_left_csr_writedata                               : out std_logic_vector(31 downto 0);                     -- writedata
			dma_comm_5_left_csr_byteenable                              : out std_logic_vector(3 downto 0);                      -- byteenable
			dma_comm_5_left_descriptor_slave_write                      : out std_logic;                                         -- write
			dma_comm_5_left_descriptor_slave_writedata                  : out std_logic_vector(255 downto 0);                    -- writedata
			dma_comm_5_left_descriptor_slave_byteenable                 : out std_logic_vector(31 downto 0);                     -- byteenable
			dma_comm_5_left_descriptor_slave_waitrequest                : in  std_logic                      := 'X';             -- waitrequest
			dma_comm_5_right_csr_address                                : out std_logic_vector(2 downto 0);                      -- address
			dma_comm_5_right_csr_write                                  : out std_logic;                                         -- write
			dma_comm_5_right_csr_read                                   : out std_logic;                                         -- read
			dma_comm_5_right_csr_readdata                               : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_comm_5_right_csr_writedata                              : out std_logic_vector(31 downto 0);                     -- writedata
			dma_comm_5_right_csr_byteenable                             : out std_logic_vector(3 downto 0);                      -- byteenable
			dma_comm_5_right_descriptor_slave_write                     : out std_logic;                                         -- write
			dma_comm_5_right_descriptor_slave_writedata                 : out std_logic_vector(255 downto 0);                    -- writedata
			dma_comm_5_right_descriptor_slave_byteenable                : out std_logic_vector(31 downto 0);                     -- byteenable
			dma_comm_5_right_descriptor_slave_waitrequest               : in  std_logic                      := 'X';             -- waitrequest
			dma_comm_6_left_csr_address                                 : out std_logic_vector(2 downto 0);                      -- address
			dma_comm_6_left_csr_write                                   : out std_logic;                                         -- write
			dma_comm_6_left_csr_read                                    : out std_logic;                                         -- read
			dma_comm_6_left_csr_readdata                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_comm_6_left_csr_writedata                               : out std_logic_vector(31 downto 0);                     -- writedata
			dma_comm_6_left_csr_byteenable                              : out std_logic_vector(3 downto 0);                      -- byteenable
			dma_comm_6_left_descriptor_slave_write                      : out std_logic;                                         -- write
			dma_comm_6_left_descriptor_slave_writedata                  : out std_logic_vector(255 downto 0);                    -- writedata
			dma_comm_6_left_descriptor_slave_byteenable                 : out std_logic_vector(31 downto 0);                     -- byteenable
			dma_comm_6_left_descriptor_slave_waitrequest                : in  std_logic                      := 'X';             -- waitrequest
			dma_comm_6_right_csr_address                                : out std_logic_vector(2 downto 0);                      -- address
			dma_comm_6_right_csr_write                                  : out std_logic;                                         -- write
			dma_comm_6_right_csr_read                                   : out std_logic;                                         -- read
			dma_comm_6_right_csr_readdata                               : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_comm_6_right_csr_writedata                              : out std_logic_vector(31 downto 0);                     -- writedata
			dma_comm_6_right_csr_byteenable                             : out std_logic_vector(3 downto 0);                      -- byteenable
			dma_comm_6_right_descriptor_slave_write                     : out std_logic;                                         -- write
			dma_comm_6_right_descriptor_slave_writedata                 : out std_logic_vector(255 downto 0);                    -- writedata
			dma_comm_6_right_descriptor_slave_byteenable                : out std_logic_vector(31 downto 0);                     -- byteenable
			dma_comm_6_right_descriptor_slave_waitrequest               : in  std_logic                      := 'X';             -- waitrequest
			dma_ftdi_usb3_csr_address                                   : out std_logic_vector(2 downto 0);                      -- address
			dma_ftdi_usb3_csr_write                                     : out std_logic;                                         -- write
			dma_ftdi_usb3_csr_read                                      : out std_logic;                                         -- read
			dma_ftdi_usb3_csr_readdata                                  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_ftdi_usb3_csr_writedata                                 : out std_logic_vector(31 downto 0);                     -- writedata
			dma_ftdi_usb3_csr_byteenable                                : out std_logic_vector(3 downto 0);                      -- byteenable
			dma_ftdi_usb3_descriptor_slave_write                        : out std_logic;                                         -- write
			dma_ftdi_usb3_descriptor_slave_writedata                    : out std_logic_vector(255 downto 0);                    -- writedata
			dma_ftdi_usb3_descriptor_slave_byteenable                   : out std_logic_vector(31 downto 0);                     -- byteenable
			dma_ftdi_usb3_descriptor_slave_waitrequest                  : in  std_logic                      := 'X';             -- waitrequest
			ext_flash_uas_address                                       : out std_logic_vector(25 downto 0);                     -- address
			ext_flash_uas_write                                         : out std_logic;                                         -- write
			ext_flash_uas_read                                          : out std_logic;                                         -- read
			ext_flash_uas_readdata                                      : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- readdata
			ext_flash_uas_writedata                                     : out std_logic_vector(15 downto 0);                     -- writedata
			ext_flash_uas_burstcount                                    : out std_logic_vector(1 downto 0);                      -- burstcount
			ext_flash_uas_byteenable                                    : out std_logic_vector(1 downto 0);                      -- byteenable
			ext_flash_uas_readdatavalid                                 : in  std_logic                      := 'X';             -- readdatavalid
			ext_flash_uas_waitrequest                                   : in  std_logic                      := 'X';             -- waitrequest
			ext_flash_uas_lock                                          : out std_logic;                                         -- lock
			ext_flash_uas_debugaccess                                   : out std_logic;                                         -- debugaccess
			FTDI_USB3_0_avalon_slave_config_address                     : out std_logic_vector(7 downto 0);                      -- address
			FTDI_USB3_0_avalon_slave_config_write                       : out std_logic;                                         -- write
			FTDI_USB3_0_avalon_slave_config_read                        : out std_logic;                                         -- read
			FTDI_USB3_0_avalon_slave_config_readdata                    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			FTDI_USB3_0_avalon_slave_config_writedata                   : out std_logic_vector(31 downto 0);                     -- writedata
			FTDI_USB3_0_avalon_slave_config_byteenable                  : out std_logic_vector(3 downto 0);                      -- byteenable
			FTDI_USB3_0_avalon_slave_config_waitrequest                 : in  std_logic                      := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_address                       : out std_logic_vector(0 downto 0);                      -- address
			jtag_uart_0_avalon_jtag_slave_write                         : out std_logic;                                         -- write
			jtag_uart_0_avalon_jtag_slave_read                          : out std_logic;                                         -- read
			jtag_uart_0_avalon_jtag_slave_readdata                      : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                     : out std_logic_vector(31 downto 0);                     -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                   : in  std_logic                      := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                    : out std_logic;                                         -- chipselect
			nios2_gen2_0_debug_mem_slave_address                        : out std_logic_vector(8 downto 0);                      -- address
			nios2_gen2_0_debug_mem_slave_write                          : out std_logic;                                         -- write
			nios2_gen2_0_debug_mem_slave_read                           : out std_logic;                                         -- read
			nios2_gen2_0_debug_mem_slave_readdata                       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                      : out std_logic_vector(31 downto 0);                     -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable                     : out std_logic_vector(3 downto 0);                      -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                    : in  std_logic                      := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                    : out std_logic;                                         -- debugaccess
			onchip_memory_s1_address                                    : out std_logic_vector(17 downto 0);                     -- address
			onchip_memory_s1_write                                      : out std_logic;                                         -- write
			onchip_memory_s1_readdata                                   : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			onchip_memory_s1_writedata                                  : out std_logic_vector(31 downto 0);                     -- writedata
			onchip_memory_s1_byteenable                                 : out std_logic_vector(3 downto 0);                      -- byteenable
			onchip_memory_s1_chipselect                                 : out std_logic;                                         -- chipselect
			onchip_memory_s1_clken                                      : out std_logic;                                         -- clken
			rmap_mem_nfee_comm_1_avalon_rmap_slave_0_address            : out std_logic_vector(11 downto 0);                     -- address
			rmap_mem_nfee_comm_1_avalon_rmap_slave_0_write              : out std_logic;                                         -- write
			rmap_mem_nfee_comm_1_avalon_rmap_slave_0_read               : out std_logic;                                         -- read
			rmap_mem_nfee_comm_1_avalon_rmap_slave_0_readdata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			rmap_mem_nfee_comm_1_avalon_rmap_slave_0_writedata          : out std_logic_vector(31 downto 0);                     -- writedata
			rmap_mem_nfee_comm_1_avalon_rmap_slave_0_byteenable         : out std_logic_vector(3 downto 0);                      -- byteenable
			rmap_mem_nfee_comm_1_avalon_rmap_slave_0_waitrequest        : in  std_logic                      := 'X';             -- waitrequest
			rmap_mem_nfee_comm_2_avalon_rmap_slave_0_address            : out std_logic_vector(11 downto 0);                     -- address
			rmap_mem_nfee_comm_2_avalon_rmap_slave_0_write              : out std_logic;                                         -- write
			rmap_mem_nfee_comm_2_avalon_rmap_slave_0_read               : out std_logic;                                         -- read
			rmap_mem_nfee_comm_2_avalon_rmap_slave_0_readdata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			rmap_mem_nfee_comm_2_avalon_rmap_slave_0_writedata          : out std_logic_vector(31 downto 0);                     -- writedata
			rmap_mem_nfee_comm_2_avalon_rmap_slave_0_byteenable         : out std_logic_vector(3 downto 0);                      -- byteenable
			rmap_mem_nfee_comm_2_avalon_rmap_slave_0_waitrequest        : in  std_logic                      := 'X';             -- waitrequest
			rmap_mem_nfee_comm_3_avalon_rmap_slave_0_address            : out std_logic_vector(11 downto 0);                     -- address
			rmap_mem_nfee_comm_3_avalon_rmap_slave_0_write              : out std_logic;                                         -- write
			rmap_mem_nfee_comm_3_avalon_rmap_slave_0_read               : out std_logic;                                         -- read
			rmap_mem_nfee_comm_3_avalon_rmap_slave_0_readdata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			rmap_mem_nfee_comm_3_avalon_rmap_slave_0_writedata          : out std_logic_vector(31 downto 0);                     -- writedata
			rmap_mem_nfee_comm_3_avalon_rmap_slave_0_byteenable         : out std_logic_vector(3 downto 0);                      -- byteenable
			rmap_mem_nfee_comm_3_avalon_rmap_slave_0_waitrequest        : in  std_logic                      := 'X';             -- waitrequest
			rmap_mem_nfee_comm_4_avalon_rmap_slave_0_address            : out std_logic_vector(11 downto 0);                     -- address
			rmap_mem_nfee_comm_4_avalon_rmap_slave_0_write              : out std_logic;                                         -- write
			rmap_mem_nfee_comm_4_avalon_rmap_slave_0_read               : out std_logic;                                         -- read
			rmap_mem_nfee_comm_4_avalon_rmap_slave_0_readdata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			rmap_mem_nfee_comm_4_avalon_rmap_slave_0_writedata          : out std_logic_vector(31 downto 0);                     -- writedata
			rmap_mem_nfee_comm_4_avalon_rmap_slave_0_byteenable         : out std_logic_vector(3 downto 0);                      -- byteenable
			rmap_mem_nfee_comm_4_avalon_rmap_slave_0_waitrequest        : in  std_logic                      := 'X';             -- waitrequest
			rmap_mem_nfee_comm_5_avalon_rmap_slave_0_address            : out std_logic_vector(11 downto 0);                     -- address
			rmap_mem_nfee_comm_5_avalon_rmap_slave_0_write              : out std_logic;                                         -- write
			rmap_mem_nfee_comm_5_avalon_rmap_slave_0_read               : out std_logic;                                         -- read
			rmap_mem_nfee_comm_5_avalon_rmap_slave_0_readdata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			rmap_mem_nfee_comm_5_avalon_rmap_slave_0_writedata          : out std_logic_vector(31 downto 0);                     -- writedata
			rmap_mem_nfee_comm_5_avalon_rmap_slave_0_byteenable         : out std_logic_vector(3 downto 0);                      -- byteenable
			rmap_mem_nfee_comm_5_avalon_rmap_slave_0_waitrequest        : in  std_logic                      := 'X';             -- waitrequest
			rmap_mem_nfee_comm_6_avalon_rmap_slave_0_address            : out std_logic_vector(11 downto 0);                     -- address
			rmap_mem_nfee_comm_6_avalon_rmap_slave_0_write              : out std_logic;                                         -- write
			rmap_mem_nfee_comm_6_avalon_rmap_slave_0_read               : out std_logic;                                         -- read
			rmap_mem_nfee_comm_6_avalon_rmap_slave_0_readdata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			rmap_mem_nfee_comm_6_avalon_rmap_slave_0_writedata          : out std_logic_vector(31 downto 0);                     -- writedata
			rmap_mem_nfee_comm_6_avalon_rmap_slave_0_byteenable         : out std_logic_vector(3 downto 0);                      -- byteenable
			rmap_mem_nfee_comm_6_avalon_rmap_slave_0_waitrequest        : in  std_logic                      := 'X';             -- waitrequest
			sysid_qsys_control_slave_address                            : out std_logic_vector(0 downto 0);                      -- address
			sysid_qsys_control_slave_readdata                           : in  std_logic_vector(31 downto 0)  := (others => 'X')  -- readdata
		);
	end component MebX_Qsys_Project_mm_interconnect_1;

	component MebX_Qsys_Project_mm_interconnect_2 is
		port (
			clk_50_clk_clk                                                         : in  std_logic                     := 'X';             -- clk
			Altera_UP_SD_Card_Avalon_Interface_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			clock_bridge_afi_50_m0_reset_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			rs232_uart_reset_reset_bridge_in_reset_reset                           : in  std_logic                     := 'X';             -- reset
			sync_reset_reset_bridge_in_reset_reset                                 : in  std_logic                     := 'X';             -- reset
			clock_bridge_afi_50_m0_address                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clock_bridge_afi_50_m0_waitrequest                                     : out std_logic;                                        -- waitrequest
			clock_bridge_afi_50_m0_burstcount                                      : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			clock_bridge_afi_50_m0_byteenable                                      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clock_bridge_afi_50_m0_read                                            : in  std_logic                     := 'X';             -- read
			clock_bridge_afi_50_m0_readdata                                        : out std_logic_vector(31 downto 0);                    -- readdata
			clock_bridge_afi_50_m0_readdatavalid                                   : out std_logic;                                        -- readdatavalid
			clock_bridge_afi_50_m0_write                                           : in  std_logic                     := 'X';             -- write
			clock_bridge_afi_50_m0_writedata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			clock_bridge_afi_50_m0_debugaccess                                     : in  std_logic                     := 'X';             -- debugaccess
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address       : out std_logic_vector(7 downto 0);                     -- address
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write         : out std_logic;                                        -- write
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read          : out std_logic;                                        -- read
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect    : out std_logic;                                        -- chipselect
			csense_adc_fo_s1_address                                               : out std_logic_vector(1 downto 0);                     -- address
			csense_adc_fo_s1_write                                                 : out std_logic;                                        -- write
			csense_adc_fo_s1_readdata                                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			csense_adc_fo_s1_writedata                                             : out std_logic_vector(31 downto 0);                    -- writedata
			csense_adc_fo_s1_chipselect                                            : out std_logic;                                        -- chipselect
			csense_cs_n_s1_address                                                 : out std_logic_vector(1 downto 0);                     -- address
			csense_cs_n_s1_write                                                   : out std_logic;                                        -- write
			csense_cs_n_s1_readdata                                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			csense_cs_n_s1_writedata                                               : out std_logic_vector(31 downto 0);                    -- writedata
			csense_cs_n_s1_chipselect                                              : out std_logic;                                        -- chipselect
			csense_sck_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			csense_sck_s1_write                                                    : out std_logic;                                        -- write
			csense_sck_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			csense_sck_s1_writedata                                                : out std_logic_vector(31 downto 0);                    -- writedata
			csense_sck_s1_chipselect                                               : out std_logic;                                        -- chipselect
			csense_sdi_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			csense_sdi_s1_write                                                    : out std_logic;                                        -- write
			csense_sdi_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			csense_sdi_s1_writedata                                                : out std_logic_vector(31 downto 0);                    -- writedata
			csense_sdi_s1_chipselect                                               : out std_logic;                                        -- chipselect
			csense_sdo_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			csense_sdo_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m1_ddr2_i2c_scl_s1_address                                             : out std_logic_vector(1 downto 0);                     -- address
			m1_ddr2_i2c_scl_s1_write                                               : out std_logic;                                        -- write
			m1_ddr2_i2c_scl_s1_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m1_ddr2_i2c_scl_s1_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			m1_ddr2_i2c_scl_s1_chipselect                                          : out std_logic;                                        -- chipselect
			m1_ddr2_i2c_sda_s1_address                                             : out std_logic_vector(1 downto 0);                     -- address
			m1_ddr2_i2c_sda_s1_write                                               : out std_logic;                                        -- write
			m1_ddr2_i2c_sda_s1_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m1_ddr2_i2c_sda_s1_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			m1_ddr2_i2c_sda_s1_chipselect                                          : out std_logic;                                        -- chipselect
			m2_ddr2_i2c_scl_s1_address                                             : out std_logic_vector(1 downto 0);                     -- address
			m2_ddr2_i2c_scl_s1_write                                               : out std_logic;                                        -- write
			m2_ddr2_i2c_scl_s1_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m2_ddr2_i2c_scl_s1_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			m2_ddr2_i2c_scl_s1_chipselect                                          : out std_logic;                                        -- chipselect
			m2_ddr2_i2c_sda_s1_address                                             : out std_logic_vector(1 downto 0);                     -- address
			m2_ddr2_i2c_sda_s1_write                                               : out std_logic;                                        -- write
			m2_ddr2_i2c_sda_s1_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m2_ddr2_i2c_sda_s1_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			m2_ddr2_i2c_sda_s1_chipselect                                          : out std_logic;                                        -- chipselect
			pio_BUTTON_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			pio_BUTTON_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_ctrl_io_lvds_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			pio_ctrl_io_lvds_s1_write                                              : out std_logic;                                        -- write
			pio_ctrl_io_lvds_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_ctrl_io_lvds_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			pio_ctrl_io_lvds_s1_chipselect                                         : out std_logic;                                        -- chipselect
			pio_DIP_s1_address                                                     : out std_logic_vector(1 downto 0);                     -- address
			pio_DIP_s1_readdata                                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_EXT_s1_address                                                     : out std_logic_vector(1 downto 0);                     -- address
			pio_EXT_s1_readdata                                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_LED_s1_address                                                     : out std_logic_vector(1 downto 0);                     -- address
			pio_LED_s1_write                                                       : out std_logic;                                        -- write
			pio_LED_s1_readdata                                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_LED_s1_writedata                                                   : out std_logic_vector(31 downto 0);                    -- writedata
			pio_LED_s1_chipselect                                                  : out std_logic;                                        -- chipselect
			pio_LED_painel_s1_address                                              : out std_logic_vector(1 downto 0);                     -- address
			pio_LED_painel_s1_write                                                : out std_logic;                                        -- write
			pio_LED_painel_s1_readdata                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_LED_painel_s1_writedata                                            : out std_logic_vector(31 downto 0);                    -- writedata
			pio_LED_painel_s1_chipselect                                           : out std_logic;                                        -- chipselect
			rs232_uart_s1_address                                                  : out std_logic_vector(2 downto 0);                     -- address
			rs232_uart_s1_write                                                    : out std_logic;                                        -- write
			rs232_uart_s1_read                                                     : out std_logic;                                        -- read
			rs232_uart_s1_readdata                                                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			rs232_uart_s1_writedata                                                : out std_logic_vector(15 downto 0);                    -- writedata
			rs232_uart_s1_begintransfer                                            : out std_logic;                                        -- begintransfer
			rs232_uart_s1_chipselect                                               : out std_logic;                                        -- chipselect
			rst_controller_avalon_rst_controller_slave_address                     : out std_logic_vector(3 downto 0);                     -- address
			rst_controller_avalon_rst_controller_slave_write                       : out std_logic;                                        -- write
			rst_controller_avalon_rst_controller_slave_read                        : out std_logic;                                        -- read
			rst_controller_avalon_rst_controller_slave_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rst_controller_avalon_rst_controller_slave_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			rst_controller_avalon_rst_controller_slave_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			rtcc_alarm_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			rtcc_alarm_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rtcc_cs_n_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			rtcc_cs_n_s1_write                                                     : out std_logic;                                        -- write
			rtcc_cs_n_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rtcc_cs_n_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			rtcc_cs_n_s1_chipselect                                                : out std_logic;                                        -- chipselect
			rtcc_sck_s1_address                                                    : out std_logic_vector(1 downto 0);                     -- address
			rtcc_sck_s1_write                                                      : out std_logic;                                        -- write
			rtcc_sck_s1_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rtcc_sck_s1_writedata                                                  : out std_logic_vector(31 downto 0);                    -- writedata
			rtcc_sck_s1_chipselect                                                 : out std_logic;                                        -- chipselect
			rtcc_sdi_s1_address                                                    : out std_logic_vector(1 downto 0);                     -- address
			rtcc_sdi_s1_write                                                      : out std_logic;                                        -- write
			rtcc_sdi_s1_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rtcc_sdi_s1_writedata                                                  : out std_logic_vector(31 downto 0);                    -- writedata
			rtcc_sdi_s1_chipselect                                                 : out std_logic;                                        -- chipselect
			rtcc_sdo_s1_address                                                    : out std_logic_vector(1 downto 0);                     -- address
			rtcc_sdo_s1_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sd_card_wp_n_s1_address                                                : out std_logic_vector(1 downto 0);                     -- address
			sd_card_wp_n_s1_readdata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SEVEN_SEGMENT_CONTROLLER_0_SSDP_avalon_slave_address                   : out std_logic_vector(0 downto 0);                     -- address
			SEVEN_SEGMENT_CONTROLLER_0_SSDP_avalon_slave_write                     : out std_logic;                                        -- write
			SEVEN_SEGMENT_CONTROLLER_0_SSDP_avalon_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			sync_avalon_mm_slave_address                                           : out std_logic_vector(7 downto 0);                     -- address
			sync_avalon_mm_slave_write                                             : out std_logic;                                        -- write
			sync_avalon_mm_slave_read                                              : out std_logic;                                        -- read
			sync_avalon_mm_slave_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sync_avalon_mm_slave_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			sync_avalon_mm_slave_byteenable                                        : out std_logic_vector(3 downto 0);                     -- byteenable
			sync_avalon_mm_slave_waitrequest                                       : in  std_logic                     := 'X';             -- waitrequest
			temp_scl_s1_address                                                    : out std_logic_vector(1 downto 0);                     -- address
			temp_scl_s1_write                                                      : out std_logic;                                        -- write
			temp_scl_s1_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			temp_scl_s1_writedata                                                  : out std_logic_vector(31 downto 0);                    -- writedata
			temp_scl_s1_chipselect                                                 : out std_logic;                                        -- chipselect
			temp_sda_s1_address                                                    : out std_logic_vector(1 downto 0);                     -- address
			temp_sda_s1_write                                                      : out std_logic;                                        -- write
			temp_sda_s1_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			temp_sda_s1_writedata                                                  : out std_logic_vector(31 downto 0);                    -- writedata
			temp_sda_s1_chipselect                                                 : out std_logic;                                        -- chipselect
			timer_1ms_s1_address                                                   : out std_logic_vector(2 downto 0);                     -- address
			timer_1ms_s1_write                                                     : out std_logic;                                        -- write
			timer_1ms_s1_readdata                                                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_1ms_s1_writedata                                                 : out std_logic_vector(15 downto 0);                    -- writedata
			timer_1ms_s1_chipselect                                                : out std_logic;                                        -- chipselect
			timer_1us_s1_address                                                   : out std_logic_vector(2 downto 0);                     -- address
			timer_1us_s1_write                                                     : out std_logic;                                        -- write
			timer_1us_s1_readdata                                                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_1us_s1_writedata                                                 : out std_logic_vector(15 downto 0);                    -- writedata
			timer_1us_s1_chipselect                                                : out std_logic                                         -- chipselect
		);
	end component MebX_Qsys_Project_mm_interconnect_2;

	component MebX_Qsys_Project_mm_interconnect_3 is
		port (
			m1_ddr2_memory_afi_clk_clk                                      : in  std_logic                      := 'X';             -- clk
			m1_ddr2_memory_afi_half_clk_clk                                 : in  std_logic                      := 'X';             -- clk
			m1_clock_bridge_m0_reset_reset_bridge_in_reset_reset            : in  std_logic                      := 'X';             -- reset
			m1_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			m1_ddr2_memory_soft_reset_reset_bridge_in_reset_reset           : in  std_logic                      := 'X';             -- reset
			m1_clock_bridge_m0_address                                      : in  std_logic_vector(30 downto 0)  := (others => 'X'); -- address
			m1_clock_bridge_m0_waitrequest                                  : out std_logic;                                         -- waitrequest
			m1_clock_bridge_m0_burstcount                                   : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- burstcount
			m1_clock_bridge_m0_byteenable                                   : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			m1_clock_bridge_m0_read                                         : in  std_logic                      := 'X';             -- read
			m1_clock_bridge_m0_readdata                                     : out std_logic_vector(255 downto 0);                    -- readdata
			m1_clock_bridge_m0_readdatavalid                                : out std_logic;                                         -- readdatavalid
			m1_clock_bridge_m0_write                                        : in  std_logic                      := 'X';             -- write
			m1_clock_bridge_m0_writedata                                    : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			m1_clock_bridge_m0_debugaccess                                  : in  std_logic                      := 'X';             -- debugaccess
			m1_ddr2_memory_avl_address                                      : out std_logic_vector(25 downto 0);                     -- address
			m1_ddr2_memory_avl_write                                        : out std_logic;                                         -- write
			m1_ddr2_memory_avl_read                                         : out std_logic;                                         -- read
			m1_ddr2_memory_avl_readdata                                     : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			m1_ddr2_memory_avl_writedata                                    : out std_logic_vector(255 downto 0);                    -- writedata
			m1_ddr2_memory_avl_beginbursttransfer                           : out std_logic;                                         -- beginbursttransfer
			m1_ddr2_memory_avl_burstcount                                   : out std_logic_vector(7 downto 0);                      -- burstcount
			m1_ddr2_memory_avl_byteenable                                   : out std_logic_vector(31 downto 0);                     -- byteenable
			m1_ddr2_memory_avl_readdatavalid                                : in  std_logic                      := 'X';             -- readdatavalid
			m1_ddr2_memory_avl_waitrequest                                  : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_3;

	component MebX_Qsys_Project_mm_interconnect_4 is
		port (
			clk_100_clk_clk                                   : in  std_logic                      := 'X';             -- clk
			dma_ftdi_usb3_reset_n_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			dma_ftdi_usb3_mm_read_address                     : in  std_logic_vector(33 downto 0)  := (others => 'X'); -- address
			dma_ftdi_usb3_mm_read_waitrequest                 : out std_logic;                                         -- waitrequest
			dma_ftdi_usb3_mm_read_byteenable                  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_ftdi_usb3_mm_read_read                        : in  std_logic                      := 'X';             -- read
			dma_ftdi_usb3_mm_read_readdata                    : out std_logic_vector(255 downto 0);                    -- readdata
			dma_ftdi_usb3_mm_read_readdatavalid               : out std_logic;                                         -- readdatavalid
			FTDI_USB3_0_avalon_slave_data_address             : out std_logic_vector(20 downto 0);                     -- address
			FTDI_USB3_0_avalon_slave_data_write               : out std_logic;                                         -- write
			FTDI_USB3_0_avalon_slave_data_read                : out std_logic;                                         -- read
			FTDI_USB3_0_avalon_slave_data_readdata            : in  std_logic_vector(255 downto 0) := (others => 'X'); -- readdata
			FTDI_USB3_0_avalon_slave_data_writedata           : out std_logic_vector(255 downto 0);                    -- writedata
			FTDI_USB3_0_avalon_slave_data_waitrequest         : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_4;

	component MebX_Qsys_Project_mm_interconnect_5 is
		port (
			clk_100_clk_clk                                              : in  std_logic                      := 'X';             -- clk
			COMM_Pedreiro_v1_01_A_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			dma_comm_1_left_reset_n_reset_bridge_in_reset_reset          : in  std_logic                      := 'X';             -- reset
			dma_comm_1_left_mm_write_address                             : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- address
			dma_comm_1_left_mm_write_waitrequest                         : out std_logic;                                         -- waitrequest
			dma_comm_1_left_mm_write_byteenable                          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_1_left_mm_write_write                               : in  std_logic                      := 'X';             -- write
			dma_comm_1_left_mm_write_writedata                           : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			COMM_Pedreiro_v1_01_A_avalon_slave_L_buffer_address          : out std_logic_vector(20 downto 0);                     -- address
			COMM_Pedreiro_v1_01_A_avalon_slave_L_buffer_write            : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_A_avalon_slave_L_buffer_writedata        : out std_logic_vector(255 downto 0);                    -- writedata
			COMM_Pedreiro_v1_01_A_avalon_slave_L_buffer_waitrequest      : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_5;

	component MebX_Qsys_Project_mm_interconnect_6 is
		port (
			clk_100_clk_clk                                              : in  std_logic                      := 'X';             -- clk
			COMM_Pedreiro_v1_01_B_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			dma_comm_2_left_reset_n_reset_bridge_in_reset_reset          : in  std_logic                      := 'X';             -- reset
			dma_comm_2_left_mm_write_address                             : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- address
			dma_comm_2_left_mm_write_waitrequest                         : out std_logic;                                         -- waitrequest
			dma_comm_2_left_mm_write_byteenable                          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_2_left_mm_write_write                               : in  std_logic                      := 'X';             -- write
			dma_comm_2_left_mm_write_writedata                           : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			COMM_Pedreiro_v1_01_B_avalon_slave_L_buffer_address          : out std_logic_vector(20 downto 0);                     -- address
			COMM_Pedreiro_v1_01_B_avalon_slave_L_buffer_write            : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_B_avalon_slave_L_buffer_writedata        : out std_logic_vector(255 downto 0);                    -- writedata
			COMM_Pedreiro_v1_01_B_avalon_slave_L_buffer_waitrequest      : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_6;

	component MebX_Qsys_Project_mm_interconnect_7 is
		port (
			clk_100_clk_clk                                              : in  std_logic                      := 'X';             -- clk
			COMM_Pedreiro_v1_01_C_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			dma_comm_3_left_reset_n_reset_bridge_in_reset_reset          : in  std_logic                      := 'X';             -- reset
			dma_comm_3_left_mm_write_address                             : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- address
			dma_comm_3_left_mm_write_waitrequest                         : out std_logic;                                         -- waitrequest
			dma_comm_3_left_mm_write_byteenable                          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_3_left_mm_write_write                               : in  std_logic                      := 'X';             -- write
			dma_comm_3_left_mm_write_writedata                           : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			COMM_Pedreiro_v1_01_C_avalon_slave_L_buffer_address          : out std_logic_vector(20 downto 0);                     -- address
			COMM_Pedreiro_v1_01_C_avalon_slave_L_buffer_write            : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_C_avalon_slave_L_buffer_writedata        : out std_logic_vector(255 downto 0);                    -- writedata
			COMM_Pedreiro_v1_01_C_avalon_slave_L_buffer_waitrequest      : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_7;

	component MebX_Qsys_Project_mm_interconnect_8 is
		port (
			clk_100_clk_clk                                              : in  std_logic                      := 'X';             -- clk
			COMM_Pedreiro_v1_01_D_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			dma_comm_4_left_reset_n_reset_bridge_in_reset_reset          : in  std_logic                      := 'X';             -- reset
			dma_comm_4_left_mm_write_address                             : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- address
			dma_comm_4_left_mm_write_waitrequest                         : out std_logic;                                         -- waitrequest
			dma_comm_4_left_mm_write_byteenable                          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_4_left_mm_write_write                               : in  std_logic                      := 'X';             -- write
			dma_comm_4_left_mm_write_writedata                           : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			COMM_Pedreiro_v1_01_D_avalon_slave_L_buffer_address          : out std_logic_vector(20 downto 0);                     -- address
			COMM_Pedreiro_v1_01_D_avalon_slave_L_buffer_write            : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_D_avalon_slave_L_buffer_writedata        : out std_logic_vector(255 downto 0);                    -- writedata
			COMM_Pedreiro_v1_01_D_avalon_slave_L_buffer_waitrequest      : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_8;

	component MebX_Qsys_Project_mm_interconnect_9 is
		port (
			clk_100_clk_clk                                              : in  std_logic                      := 'X';             -- clk
			COMM_Pedreiro_v1_01_E_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			dma_comm_5_left_reset_n_reset_bridge_in_reset_reset          : in  std_logic                      := 'X';             -- reset
			dma_comm_5_left_mm_write_address                             : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- address
			dma_comm_5_left_mm_write_waitrequest                         : out std_logic;                                         -- waitrequest
			dma_comm_5_left_mm_write_byteenable                          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_5_left_mm_write_write                               : in  std_logic                      := 'X';             -- write
			dma_comm_5_left_mm_write_writedata                           : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			COMM_Pedreiro_v1_01_E_avalon_slave_L_buffer_address          : out std_logic_vector(20 downto 0);                     -- address
			COMM_Pedreiro_v1_01_E_avalon_slave_L_buffer_write            : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_E_avalon_slave_L_buffer_writedata        : out std_logic_vector(255 downto 0);                    -- writedata
			COMM_Pedreiro_v1_01_E_avalon_slave_L_buffer_waitrequest      : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_9;

	component MebX_Qsys_Project_mm_interconnect_10 is
		port (
			clk_100_clk_clk                                              : in  std_logic                      := 'X';             -- clk
			COMM_Pedreiro_v1_01_F_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			dma_comm_6_left_reset_n_reset_bridge_in_reset_reset          : in  std_logic                      := 'X';             -- reset
			dma_comm_6_left_mm_write_address                             : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- address
			dma_comm_6_left_mm_write_waitrequest                         : out std_logic;                                         -- waitrequest
			dma_comm_6_left_mm_write_byteenable                          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_6_left_mm_write_write                               : in  std_logic                      := 'X';             -- write
			dma_comm_6_left_mm_write_writedata                           : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			COMM_Pedreiro_v1_01_F_avalon_slave_L_buffer_address          : out std_logic_vector(20 downto 0);                     -- address
			COMM_Pedreiro_v1_01_F_avalon_slave_L_buffer_write            : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_F_avalon_slave_L_buffer_writedata        : out std_logic_vector(255 downto 0);                    -- writedata
			COMM_Pedreiro_v1_01_F_avalon_slave_L_buffer_waitrequest      : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_10;

	component MebX_Qsys_Project_mm_interconnect_11 is
		port (
			clk_100_clk_clk                                              : in  std_logic                      := 'X';             -- clk
			COMM_Pedreiro_v1_01_A_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			dma_comm_1_right_reset_n_reset_bridge_in_reset_reset         : in  std_logic                      := 'X';             -- reset
			dma_comm_1_right_mm_write_address                            : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- address
			dma_comm_1_right_mm_write_waitrequest                        : out std_logic;                                         -- waitrequest
			dma_comm_1_right_mm_write_byteenable                         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_1_right_mm_write_write                              : in  std_logic                      := 'X';             -- write
			dma_comm_1_right_mm_write_writedata                          : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			COMM_Pedreiro_v1_01_A_avalon_slave_R_buffer_address          : out std_logic_vector(20 downto 0);                     -- address
			COMM_Pedreiro_v1_01_A_avalon_slave_R_buffer_write            : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_A_avalon_slave_R_buffer_writedata        : out std_logic_vector(255 downto 0);                    -- writedata
			COMM_Pedreiro_v1_01_A_avalon_slave_R_buffer_waitrequest      : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_11;

	component MebX_Qsys_Project_mm_interconnect_12 is
		port (
			clk_100_clk_clk                                              : in  std_logic                      := 'X';             -- clk
			COMM_Pedreiro_v1_01_B_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			dma_comm_2_right_reset_n_reset_bridge_in_reset_reset         : in  std_logic                      := 'X';             -- reset
			dma_comm_2_right_mm_write_address                            : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- address
			dma_comm_2_right_mm_write_waitrequest                        : out std_logic;                                         -- waitrequest
			dma_comm_2_right_mm_write_byteenable                         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_2_right_mm_write_write                              : in  std_logic                      := 'X';             -- write
			dma_comm_2_right_mm_write_writedata                          : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			COMM_Pedreiro_v1_01_B_avalon_slave_R_buffer_address          : out std_logic_vector(20 downto 0);                     -- address
			COMM_Pedreiro_v1_01_B_avalon_slave_R_buffer_write            : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_B_avalon_slave_R_buffer_writedata        : out std_logic_vector(255 downto 0);                    -- writedata
			COMM_Pedreiro_v1_01_B_avalon_slave_R_buffer_waitrequest      : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_12;

	component MebX_Qsys_Project_mm_interconnect_13 is
		port (
			clk_100_clk_clk                                              : in  std_logic                      := 'X';             -- clk
			COMM_Pedreiro_v1_01_C_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			dma_comm_3_right_reset_n_reset_bridge_in_reset_reset         : in  std_logic                      := 'X';             -- reset
			dma_comm_3_right_mm_write_address                            : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- address
			dma_comm_3_right_mm_write_waitrequest                        : out std_logic;                                         -- waitrequest
			dma_comm_3_right_mm_write_byteenable                         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_3_right_mm_write_write                              : in  std_logic                      := 'X';             -- write
			dma_comm_3_right_mm_write_writedata                          : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			COMM_Pedreiro_v1_01_C_avalon_slave_R_buffer_address          : out std_logic_vector(20 downto 0);                     -- address
			COMM_Pedreiro_v1_01_C_avalon_slave_R_buffer_write            : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_C_avalon_slave_R_buffer_writedata        : out std_logic_vector(255 downto 0);                    -- writedata
			COMM_Pedreiro_v1_01_C_avalon_slave_R_buffer_waitrequest      : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_13;

	component MebX_Qsys_Project_mm_interconnect_14 is
		port (
			clk_100_clk_clk                                              : in  std_logic                      := 'X';             -- clk
			COMM_Pedreiro_v1_01_D_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			dma_comm_4_right_reset_n_reset_bridge_in_reset_reset         : in  std_logic                      := 'X';             -- reset
			dma_comm_4_right_mm_write_address                            : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- address
			dma_comm_4_right_mm_write_waitrequest                        : out std_logic;                                         -- waitrequest
			dma_comm_4_right_mm_write_byteenable                         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_4_right_mm_write_write                              : in  std_logic                      := 'X';             -- write
			dma_comm_4_right_mm_write_writedata                          : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			COMM_Pedreiro_v1_01_D_avalon_slave_R_buffer_address          : out std_logic_vector(20 downto 0);                     -- address
			COMM_Pedreiro_v1_01_D_avalon_slave_R_buffer_write            : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_D_avalon_slave_R_buffer_writedata        : out std_logic_vector(255 downto 0);                    -- writedata
			COMM_Pedreiro_v1_01_D_avalon_slave_R_buffer_waitrequest      : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_14;

	component MebX_Qsys_Project_mm_interconnect_15 is
		port (
			clk_100_clk_clk                                              : in  std_logic                      := 'X';             -- clk
			COMM_Pedreiro_v1_01_E_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			dma_comm_5_right_reset_n_reset_bridge_in_reset_reset         : in  std_logic                      := 'X';             -- reset
			dma_comm_5_right_mm_write_address                            : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- address
			dma_comm_5_right_mm_write_waitrequest                        : out std_logic;                                         -- waitrequest
			dma_comm_5_right_mm_write_byteenable                         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_5_right_mm_write_write                              : in  std_logic                      := 'X';             -- write
			dma_comm_5_right_mm_write_writedata                          : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			COMM_Pedreiro_v1_01_E_avalon_slave_R_buffer_address          : out std_logic_vector(20 downto 0);                     -- address
			COMM_Pedreiro_v1_01_E_avalon_slave_R_buffer_write            : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_E_avalon_slave_R_buffer_writedata        : out std_logic_vector(255 downto 0);                    -- writedata
			COMM_Pedreiro_v1_01_E_avalon_slave_R_buffer_waitrequest      : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_15;

	component MebX_Qsys_Project_mm_interconnect_16 is
		port (
			clk_100_clk_clk                                              : in  std_logic                      := 'X';             -- clk
			COMM_Pedreiro_v1_01_F_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			dma_comm_6_right_reset_n_reset_bridge_in_reset_reset         : in  std_logic                      := 'X';             -- reset
			dma_comm_6_right_mm_write_address                            : in  std_logic_vector(32 downto 0)  := (others => 'X'); -- address
			dma_comm_6_right_mm_write_waitrequest                        : out std_logic;                                         -- waitrequest
			dma_comm_6_right_mm_write_byteenable                         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			dma_comm_6_right_mm_write_write                              : in  std_logic                      := 'X';             -- write
			dma_comm_6_right_mm_write_writedata                          : in  std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			COMM_Pedreiro_v1_01_F_avalon_slave_R_buffer_address          : out std_logic_vector(20 downto 0);                     -- address
			COMM_Pedreiro_v1_01_F_avalon_slave_R_buffer_write            : out std_logic;                                         -- write
			COMM_Pedreiro_v1_01_F_avalon_slave_R_buffer_writedata        : out std_logic_vector(255 downto 0);                    -- writedata
			COMM_Pedreiro_v1_01_F_avalon_slave_R_buffer_waitrequest      : in  std_logic                      := 'X'              -- waitrequest
		);
	end component MebX_Qsys_Project_mm_interconnect_16;

	component MebX_Qsys_Project_irq_mapper is
		port (
			clk            : in  std_logic                     := 'X'; -- clk
			reset          : in  std_logic                     := 'X'; -- reset
			receiver0_irq  : in  std_logic                     := 'X'; -- irq
			receiver1_irq  : in  std_logic                     := 'X'; -- irq
			receiver2_irq  : in  std_logic                     := 'X'; -- irq
			receiver3_irq  : in  std_logic                     := 'X'; -- irq
			receiver4_irq  : in  std_logic                     := 'X'; -- irq
			receiver5_irq  : in  std_logic                     := 'X'; -- irq
			receiver6_irq  : in  std_logic                     := 'X'; -- irq
			receiver7_irq  : in  std_logic                     := 'X'; -- irq
			receiver8_irq  : in  std_logic                     := 'X'; -- irq
			receiver9_irq  : in  std_logic                     := 'X'; -- irq
			receiver10_irq : in  std_logic                     := 'X'; -- irq
			receiver11_irq : in  std_logic                     := 'X'; -- irq
			receiver12_irq : in  std_logic                     := 'X'; -- irq
			receiver13_irq : in  std_logic                     := 'X'; -- irq
			receiver14_irq : in  std_logic                     := 'X'; -- irq
			receiver15_irq : in  std_logic                     := 'X'; -- irq
			receiver16_irq : in  std_logic                     := 'X'; -- irq
			receiver17_irq : in  std_logic                     := 'X'; -- irq
			receiver18_irq : in  std_logic                     := 'X'; -- irq
			receiver19_irq : in  std_logic                     := 'X'; -- irq
			receiver20_irq : in  std_logic                     := 'X'; -- irq
			receiver21_irq : in  std_logic                     := 'X'; -- irq
			receiver22_irq : in  std_logic                     := 'X'; -- irq
			receiver23_irq : in  std_logic                     := 'X'; -- irq
			receiver24_irq : in  std_logic                     := 'X'; -- irq
			receiver25_irq : in  std_logic                     := 'X'; -- irq
			receiver26_irq : in  std_logic                     := 'X'; -- irq
			receiver27_irq : in  std_logic                     := 'X'; -- irq
			receiver28_irq : in  std_logic                     := 'X'; -- irq
			receiver29_irq : in  std_logic                     := 'X'; -- irq
			receiver30_irq : in  std_logic                     := 'X'; -- irq
			receiver31_irq : in  std_logic                     := 'X'; -- irq
			sender_irq     : out std_logic_vector(31 downto 0)         -- irq
		);
	end component MebX_Qsys_Project_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component mebx_qsys_project_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component mebx_qsys_project_rst_controller_001;

	component mebx_qsys_project_rst_controller_008 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component mebx_qsys_project_rst_controller_008;

	component mebx_qsys_project_rst_controller_009 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component mebx_qsys_project_rst_controller_009;

	component mebx_qsys_project_clock_bridge_afi_50 is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			HDL_ADDR_WIDTH      : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             --   m0_clk.clk
			m0_reset         : in  std_logic                     := 'X';             -- m0_reset.reset
			s0_clk           : in  std_logic                     := 'X';             --   s0_clk.clk
			s0_reset         : in  std_logic                     := 'X';             -- s0_reset.reset
			s0_waitrequest   : out std_logic;                                        --       s0.waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    --         .readdata
			s0_readdatavalid : out std_logic;                                        --         .readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); --         .burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); --         .writedata
			s0_address       : in  std_logic_vector(11 downto 0) := (others => 'X'); --         .address
			s0_write         : in  std_logic                     := 'X';             --         .write
			s0_read          : in  std_logic                     := 'X';             --         .read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); --         .byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             --         .debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             --       m0.waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); --         .readdata
			m0_readdatavalid : in  std_logic                     := 'X';             --         .readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     --         .burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    --         .writedata
			m0_address       : out std_logic_vector(11 downto 0);                    --         .address
			m0_write         : out std_logic;                                        --         .write
			m0_read          : out std_logic;                                        --         .read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     --         .byteenable
			m0_debugaccess   : out std_logic                                         --         .debugaccess
		);
	end component mebx_qsys_project_clock_bridge_afi_50;

	component mebx_qsys_project_m1_clock_bridge is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			HDL_ADDR_WIDTH      : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                      := 'X';             --   m0_clk.clk
			m0_reset         : in  std_logic                      := 'X';             -- m0_reset.reset
			s0_clk           : in  std_logic                      := 'X';             --   s0_clk.clk
			s0_reset         : in  std_logic                      := 'X';             -- s0_reset.reset
			s0_waitrequest   : out std_logic;                                         --       s0.waitrequest
			s0_readdata      : out std_logic_vector(255 downto 0);                    --         .readdata
			s0_readdatavalid : out std_logic;                                         --         .readdatavalid
			s0_burstcount    : in  std_logic_vector(2 downto 0)   := (others => 'X'); --         .burstcount
			s0_writedata     : in  std_logic_vector(255 downto 0) := (others => 'X'); --         .writedata
			s0_address       : in  std_logic_vector(30 downto 0)  := (others => 'X'); --         .address
			s0_write         : in  std_logic                      := 'X';             --         .write
			s0_read          : in  std_logic                      := 'X';             --         .read
			s0_byteenable    : in  std_logic_vector(31 downto 0)  := (others => 'X'); --         .byteenable
			s0_debugaccess   : in  std_logic                      := 'X';             --         .debugaccess
			m0_waitrequest   : in  std_logic                      := 'X';             --       m0.waitrequest
			m0_readdata      : in  std_logic_vector(255 downto 0) := (others => 'X'); --         .readdata
			m0_readdatavalid : in  std_logic                      := 'X';             --         .readdatavalid
			m0_burstcount    : out std_logic_vector(2 downto 0);                      --         .burstcount
			m0_writedata     : out std_logic_vector(255 downto 0);                    --         .writedata
			m0_address       : out std_logic_vector(30 downto 0);                     --         .address
			m0_write         : out std_logic;                                         --         .write
			m0_read          : out std_logic;                                         --         .read
			m0_byteenable    : out std_logic_vector(31 downto 0);                     --         .byteenable
			m0_debugaccess   : out std_logic                                          --         .debugaccess
		);
	end component mebx_qsys_project_m1_clock_bridge;

	signal m2_ddr2_memory_afi_clk_clk                                                             : std_logic;                      -- m2_ddr2_memory:afi_clk -> [COMM_Pedreiro_v1_01_A:clock_sink_200_clk, COMM_Pedreiro_v1_01_B:clock_sink_200_clk, COMM_Pedreiro_v1_01_C:clock_sink_200_clk, COMM_Pedreiro_v1_01_D:clock_sink_200_clk, COMM_Pedreiro_v1_01_E:clock_sink_200_clk, COMM_Pedreiro_v1_01_F:clock_sink_200_clk, mm_interconnect_0:m2_ddr2_memory_afi_clk_clk, rst_controller_015:clk]
	signal m2_ddr2_memory_afi_half_clk_clk                                                        : std_logic;                      -- m2_ddr2_memory:afi_half_clk -> [COMM_Pedreiro_v1_01_A:clock_sink_100_clk, COMM_Pedreiro_v1_01_B:clock_sink_100_clk, COMM_Pedreiro_v1_01_C:clock_sink_100_clk, COMM_Pedreiro_v1_01_D:clock_sink_100_clk, COMM_Pedreiro_v1_01_E:clock_sink_100_clk, COMM_Pedreiro_v1_01_F:clock_sink_100_clk, FTDI_USB3_0:clock_sink_clk, clock_bridge_afi_50:s0_clk, ddr2_address_span_extender:clk, dma_comm_1_left:clock_clk, dma_comm_1_right:clock_clk, dma_comm_2_left:clock_clk, dma_comm_2_right:clock_clk, dma_comm_3_left:clock_clk, dma_comm_3_right:clock_clk, dma_comm_4_left:clock_clk, dma_comm_4_right:clock_clk, dma_comm_5_left:clock_clk, dma_comm_5_right:clock_clk, dma_comm_6_left:clock_clk, dma_comm_6_right:clock_clk, dma_ftdi_usb3:clock_clk, ext_flash:clk_clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, irq_synchronizer_004:sender_clk, jtag_uart_0:clk, m1_clock_bridge:s0_clk, mm_interconnect_0:clk_100_clk_clk, mm_interconnect_0:m2_ddr2_memory_afi_half_clk_clk, mm_interconnect_10:clk_100_clk_clk, mm_interconnect_11:clk_100_clk_clk, mm_interconnect_12:clk_100_clk_clk, mm_interconnect_13:clk_100_clk_clk, mm_interconnect_14:clk_100_clk_clk, mm_interconnect_15:clk_100_clk_clk, mm_interconnect_16:clk_100_clk_clk, mm_interconnect_1:clk_100_clk_clk, mm_interconnect_4:clk_100_clk_clk, mm_interconnect_5:clk_100_clk_clk, mm_interconnect_6:clk_100_clk_clk, mm_interconnect_7:clk_100_clk_clk, mm_interconnect_8:clk_100_clk_clk, mm_interconnect_9:clk_100_clk_clk, nios2_gen2_0:clk, onchip_memory:clk, rmap_mem_nfee_comm_1:clk_100_i, rmap_mem_nfee_comm_2:clk_100_i, rmap_mem_nfee_comm_3:clk_100_i, rmap_mem_nfee_comm_4:clk_100_i, rmap_mem_nfee_comm_5:clk_100_i, rmap_mem_nfee_comm_6:clk_100_i, rst_controller_002:clk, rst_controller_003:clk, rst_controller_004:clk, rst_controller_005:clk, rst_controller_006:clk, rst_controller_007:clk, rst_controller_008:clk, rst_controller_010:clk, rst_controller_012:clk, sysid_qsys:clock, tristate_conduit_bridge_0:clk]
	signal m1_ddr2_memory_afi_half_clk_clk                                                        : std_logic;                      -- m1_ddr2_memory:afi_half_clk -> [m1_clock_bridge:m0_clk, mm_interconnect_3:m1_ddr2_memory_afi_half_clk_clk, rst_controller_011:clk]
	signal comm_pedreiro_v1_01_a_conduit_end_avm_configs_out_win_mem_addr_offset_signal           : std_logic_vector(63 downto 0);  -- COMM_Pedreiro_v1_01_A:channel_win_mem_addr_offset_o -> rmap_mem_nfee_comm_1:channel_win_mem_addr_offset_i
	signal comm_pedreiro_v1_01_c_conduit_end_avm_configs_out_win_mem_addr_offset_signal           : std_logic_vector(63 downto 0);  -- COMM_Pedreiro_v1_01_C:channel_win_mem_addr_offset_o -> rmap_mem_nfee_comm_3:channel_win_mem_addr_offset_i
	signal comm_pedreiro_v1_01_b_conduit_end_avm_configs_out_win_mem_addr_offset_signal           : std_logic_vector(63 downto 0);  -- COMM_Pedreiro_v1_01_B:channel_win_mem_addr_offset_o -> rmap_mem_nfee_comm_2:channel_win_mem_addr_offset_i
	signal comm_pedreiro_v1_01_d_conduit_end_avm_configs_out_win_mem_addr_offset_signal           : std_logic_vector(63 downto 0);  -- COMM_Pedreiro_v1_01_D:channel_win_mem_addr_offset_o -> rmap_mem_nfee_comm_4:channel_win_mem_addr_offset_i
	signal comm_pedreiro_v1_01_e_conduit_end_avm_configs_out_win_mem_addr_offset_signal           : std_logic_vector(63 downto 0);  -- COMM_Pedreiro_v1_01_E:channel_win_mem_addr_offset_o -> rmap_mem_nfee_comm_5:channel_win_mem_addr_offset_i
	signal comm_pedreiro_v1_01_f_conduit_end_avm_configs_out_win_mem_addr_offset_signal           : std_logic_vector(63 downto 0);  -- COMM_Pedreiro_v1_01_F:channel_win_mem_addr_offset_o -> rmap_mem_nfee_comm_6:channel_win_mem_addr_offset_i
	signal comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_timecode_time_signal                  : std_logic_vector(5 downto 0);   -- COMM_Pedreiro_v1_01_A:channel_hk_timecode_time_o -> rmap_mem_nfee_comm_1:channel_hk_timecode_time_i
	signal comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_parity_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_A:channel_hk_spw_link_parity_err_o -> rmap_mem_nfee_comm_1:channel_hk_spw_link_parity_err_i
	signal comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_disconnect_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_A:channel_hk_spw_link_disconnect_o -> rmap_mem_nfee_comm_1:channel_hk_spw_link_disconnect_i
	signal comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_escape_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_A:channel_hk_spw_link_escape_err_o -> rmap_mem_nfee_comm_1:channel_hk_spw_link_escape_err_i
	signal comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_rmap_target_indicate_signal           : std_logic;                      -- COMM_Pedreiro_v1_01_A:channel_hk_rmap_target_indicate_o -> rmap_mem_nfee_comm_1:channel_hk_rmap_target_indicate_i
	signal comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_running_signal               : std_logic;                      -- COMM_Pedreiro_v1_01_A:channel_hk_spw_link_running_o -> rmap_mem_nfee_comm_1:channel_hk_spw_link_running_i
	signal comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_frame_counter_signal                  : std_logic_vector(15 downto 0);  -- COMM_Pedreiro_v1_01_A:channel_hk_frame_counter_o -> rmap_mem_nfee_comm_1:channel_hk_frame_counter_i
	signal comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_credit_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_A:channel_hk_spw_link_credit_err_o -> rmap_mem_nfee_comm_1:channel_hk_spw_link_credit_err_i
	signal comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_timecode_control_signal               : std_logic_vector(1 downto 0);   -- COMM_Pedreiro_v1_01_A:channel_hk_timecode_control_o -> rmap_mem_nfee_comm_1:channel_hk_timecode_control_i
	signal comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_frame_number_signal                   : std_logic_vector(1 downto 0);   -- COMM_Pedreiro_v1_01_A:channel_hk_frame_number_o -> rmap_mem_nfee_comm_1:channel_hk_frame_number_i
	signal comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_rmap_target_status_signal             : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_A:channel_hk_rmap_target_status_o -> rmap_mem_nfee_comm_1:channel_hk_rmap_target_status_i
	signal comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_timecode_time_signal                  : std_logic_vector(5 downto 0);   -- COMM_Pedreiro_v1_01_B:channel_hk_timecode_time_o -> rmap_mem_nfee_comm_2:channel_hk_timecode_time_i
	signal comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_parity_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_B:channel_hk_spw_link_parity_err_o -> rmap_mem_nfee_comm_2:channel_hk_spw_link_parity_err_i
	signal comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_disconnect_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_B:channel_hk_spw_link_disconnect_o -> rmap_mem_nfee_comm_2:channel_hk_spw_link_disconnect_i
	signal comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_escape_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_B:channel_hk_spw_link_escape_err_o -> rmap_mem_nfee_comm_2:channel_hk_spw_link_escape_err_i
	signal comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_rmap_target_indicate_signal           : std_logic;                      -- COMM_Pedreiro_v1_01_B:channel_hk_rmap_target_indicate_o -> rmap_mem_nfee_comm_2:channel_hk_rmap_target_indicate_i
	signal comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_running_signal               : std_logic;                      -- COMM_Pedreiro_v1_01_B:channel_hk_spw_link_running_o -> rmap_mem_nfee_comm_2:channel_hk_spw_link_running_i
	signal comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_frame_counter_signal                  : std_logic_vector(15 downto 0);  -- COMM_Pedreiro_v1_01_B:channel_hk_frame_counter_o -> rmap_mem_nfee_comm_2:channel_hk_frame_counter_i
	signal comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_credit_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_B:channel_hk_spw_link_credit_err_o -> rmap_mem_nfee_comm_2:channel_hk_spw_link_credit_err_i
	signal comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_timecode_control_signal               : std_logic_vector(1 downto 0);   -- COMM_Pedreiro_v1_01_B:channel_hk_timecode_control_o -> rmap_mem_nfee_comm_2:channel_hk_timecode_control_i
	signal comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_frame_number_signal                   : std_logic_vector(1 downto 0);   -- COMM_Pedreiro_v1_01_B:channel_hk_frame_number_o -> rmap_mem_nfee_comm_2:channel_hk_frame_number_i
	signal comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_rmap_target_status_signal             : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_B:channel_hk_rmap_target_status_o -> rmap_mem_nfee_comm_2:channel_hk_rmap_target_status_i
	signal comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_timecode_time_signal                  : std_logic_vector(5 downto 0);   -- COMM_Pedreiro_v1_01_C:channel_hk_timecode_time_o -> rmap_mem_nfee_comm_3:channel_hk_timecode_time_i
	signal comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_parity_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_C:channel_hk_spw_link_parity_err_o -> rmap_mem_nfee_comm_3:channel_hk_spw_link_parity_err_i
	signal comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_disconnect_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_C:channel_hk_spw_link_disconnect_o -> rmap_mem_nfee_comm_3:channel_hk_spw_link_disconnect_i
	signal comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_escape_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_C:channel_hk_spw_link_escape_err_o -> rmap_mem_nfee_comm_3:channel_hk_spw_link_escape_err_i
	signal comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_rmap_target_indicate_signal           : std_logic;                      -- COMM_Pedreiro_v1_01_C:channel_hk_rmap_target_indicate_o -> rmap_mem_nfee_comm_3:channel_hk_rmap_target_indicate_i
	signal comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_running_signal               : std_logic;                      -- COMM_Pedreiro_v1_01_C:channel_hk_spw_link_running_o -> rmap_mem_nfee_comm_3:channel_hk_spw_link_running_i
	signal comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_frame_counter_signal                  : std_logic_vector(15 downto 0);  -- COMM_Pedreiro_v1_01_C:channel_hk_frame_counter_o -> rmap_mem_nfee_comm_3:channel_hk_frame_counter_i
	signal comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_credit_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_C:channel_hk_spw_link_credit_err_o -> rmap_mem_nfee_comm_3:channel_hk_spw_link_credit_err_i
	signal comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_timecode_control_signal               : std_logic_vector(1 downto 0);   -- COMM_Pedreiro_v1_01_C:channel_hk_timecode_control_o -> rmap_mem_nfee_comm_3:channel_hk_timecode_control_i
	signal comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_frame_number_signal                   : std_logic_vector(1 downto 0);   -- COMM_Pedreiro_v1_01_C:channel_hk_frame_number_o -> rmap_mem_nfee_comm_3:channel_hk_frame_number_i
	signal comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_rmap_target_status_signal             : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_C:channel_hk_rmap_target_status_o -> rmap_mem_nfee_comm_3:channel_hk_rmap_target_status_i
	signal comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_timecode_time_signal                  : std_logic_vector(5 downto 0);   -- COMM_Pedreiro_v1_01_D:channel_hk_timecode_time_o -> rmap_mem_nfee_comm_4:channel_hk_timecode_time_i
	signal comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_parity_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_D:channel_hk_spw_link_parity_err_o -> rmap_mem_nfee_comm_4:channel_hk_spw_link_parity_err_i
	signal comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_disconnect_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_D:channel_hk_spw_link_disconnect_o -> rmap_mem_nfee_comm_4:channel_hk_spw_link_disconnect_i
	signal comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_escape_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_D:channel_hk_spw_link_escape_err_o -> rmap_mem_nfee_comm_4:channel_hk_spw_link_escape_err_i
	signal comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_rmap_target_indicate_signal           : std_logic;                      -- COMM_Pedreiro_v1_01_D:channel_hk_rmap_target_indicate_o -> rmap_mem_nfee_comm_4:channel_hk_rmap_target_indicate_i
	signal comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_running_signal               : std_logic;                      -- COMM_Pedreiro_v1_01_D:channel_hk_spw_link_running_o -> rmap_mem_nfee_comm_4:channel_hk_spw_link_running_i
	signal comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_frame_counter_signal                  : std_logic_vector(15 downto 0);  -- COMM_Pedreiro_v1_01_D:channel_hk_frame_counter_o -> rmap_mem_nfee_comm_4:channel_hk_frame_counter_i
	signal comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_credit_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_D:channel_hk_spw_link_credit_err_o -> rmap_mem_nfee_comm_4:channel_hk_spw_link_credit_err_i
	signal comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_timecode_control_signal               : std_logic_vector(1 downto 0);   -- COMM_Pedreiro_v1_01_D:channel_hk_timecode_control_o -> rmap_mem_nfee_comm_4:channel_hk_timecode_control_i
	signal comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_frame_number_signal                   : std_logic_vector(1 downto 0);   -- COMM_Pedreiro_v1_01_D:channel_hk_frame_number_o -> rmap_mem_nfee_comm_4:channel_hk_frame_number_i
	signal comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_rmap_target_status_signal             : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_D:channel_hk_rmap_target_status_o -> rmap_mem_nfee_comm_4:channel_hk_rmap_target_status_i
	signal comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_timecode_time_signal                  : std_logic_vector(5 downto 0);   -- COMM_Pedreiro_v1_01_F:channel_hk_timecode_time_o -> rmap_mem_nfee_comm_6:channel_hk_timecode_time_i
	signal comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_parity_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_F:channel_hk_spw_link_parity_err_o -> rmap_mem_nfee_comm_6:channel_hk_spw_link_parity_err_i
	signal comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_disconnect_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_F:channel_hk_spw_link_disconnect_o -> rmap_mem_nfee_comm_6:channel_hk_spw_link_disconnect_i
	signal comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_escape_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_F:channel_hk_spw_link_escape_err_o -> rmap_mem_nfee_comm_6:channel_hk_spw_link_escape_err_i
	signal comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_rmap_target_indicate_signal           : std_logic;                      -- COMM_Pedreiro_v1_01_F:channel_hk_rmap_target_indicate_o -> rmap_mem_nfee_comm_6:channel_hk_rmap_target_indicate_i
	signal comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_running_signal               : std_logic;                      -- COMM_Pedreiro_v1_01_F:channel_hk_spw_link_running_o -> rmap_mem_nfee_comm_6:channel_hk_spw_link_running_i
	signal comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_frame_counter_signal                  : std_logic_vector(15 downto 0);  -- COMM_Pedreiro_v1_01_F:channel_hk_frame_counter_o -> rmap_mem_nfee_comm_6:channel_hk_frame_counter_i
	signal comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_credit_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_F:channel_hk_spw_link_credit_err_o -> rmap_mem_nfee_comm_6:channel_hk_spw_link_credit_err_i
	signal comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_timecode_control_signal               : std_logic_vector(1 downto 0);   -- COMM_Pedreiro_v1_01_F:channel_hk_timecode_control_o -> rmap_mem_nfee_comm_6:channel_hk_timecode_control_i
	signal comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_frame_number_signal                   : std_logic_vector(1 downto 0);   -- COMM_Pedreiro_v1_01_F:channel_hk_frame_number_o -> rmap_mem_nfee_comm_6:channel_hk_frame_number_i
	signal comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_rmap_target_status_signal             : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_F:channel_hk_rmap_target_status_o -> rmap_mem_nfee_comm_6:channel_hk_rmap_target_status_i
	signal comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_timecode_time_signal                  : std_logic_vector(5 downto 0);   -- COMM_Pedreiro_v1_01_E:channel_hk_timecode_time_o -> rmap_mem_nfee_comm_5:channel_hk_timecode_time_i
	signal comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_parity_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_E:channel_hk_spw_link_parity_err_o -> rmap_mem_nfee_comm_5:channel_hk_spw_link_parity_err_i
	signal comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_disconnect_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_E:channel_hk_spw_link_disconnect_o -> rmap_mem_nfee_comm_5:channel_hk_spw_link_disconnect_i
	signal comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_escape_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_E:channel_hk_spw_link_escape_err_o -> rmap_mem_nfee_comm_5:channel_hk_spw_link_escape_err_i
	signal comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_rmap_target_indicate_signal           : std_logic;                      -- COMM_Pedreiro_v1_01_E:channel_hk_rmap_target_indicate_o -> rmap_mem_nfee_comm_5:channel_hk_rmap_target_indicate_i
	signal comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_running_signal               : std_logic;                      -- COMM_Pedreiro_v1_01_E:channel_hk_spw_link_running_o -> rmap_mem_nfee_comm_5:channel_hk_spw_link_running_i
	signal comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_frame_counter_signal                  : std_logic_vector(15 downto 0);  -- COMM_Pedreiro_v1_01_E:channel_hk_frame_counter_o -> rmap_mem_nfee_comm_5:channel_hk_frame_counter_i
	signal comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_credit_err_signal            : std_logic;                      -- COMM_Pedreiro_v1_01_E:channel_hk_spw_link_credit_err_o -> rmap_mem_nfee_comm_5:channel_hk_spw_link_credit_err_i
	signal comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_timecode_control_signal               : std_logic_vector(1 downto 0);   -- COMM_Pedreiro_v1_01_E:channel_hk_timecode_control_o -> rmap_mem_nfee_comm_5:channel_hk_timecode_control_i
	signal comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_frame_number_signal                   : std_logic_vector(1 downto 0);   -- COMM_Pedreiro_v1_01_E:channel_hk_frame_number_o -> rmap_mem_nfee_comm_5:channel_hk_frame_number_i
	signal comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_rmap_target_status_signal             : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_E:channel_hk_rmap_target_status_o -> rmap_mem_nfee_comm_5:channel_hk_rmap_target_status_i
	signal comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_write_signal                   : std_logic;                      -- COMM_Pedreiro_v1_01_C:fee_codec_rmap_write_o -> rmap_mem_nfee_comm_3:fee_0_rmap_write_i
	signal rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_readdata_signal                      : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_3:fee_0_rmap_readdata_o -> COMM_Pedreiro_v1_01_C:fee_codec_rmap_readdata_i
	signal comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_rd_address_signal              : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_C:fee_codec_rmap_rd_address_o -> rmap_mem_nfee_comm_3:fee_0_rmap_rd_address_i
	signal comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_wr_address_signal              : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_C:fee_codec_rmap_wr_address_o -> rmap_mem_nfee_comm_3:fee_0_rmap_wr_address_i
	signal comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_read_signal                    : std_logic;                      -- COMM_Pedreiro_v1_01_C:fee_codec_rmap_read_o -> rmap_mem_nfee_comm_3:fee_0_rmap_read_i
	signal rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_3:fee_0_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_C:fee_codec_rmap_wr_waitrequest_i
	signal rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_3:fee_0_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_C:fee_codec_rmap_rd_waitrequest_i
	signal comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_writedata_signal               : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_C:fee_codec_rmap_writedata_o -> rmap_mem_nfee_comm_3:fee_0_rmap_writedata_i
	signal comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_write_signal                   : std_logic;                      -- COMM_Pedreiro_v1_01_A:fee_codec_rmap_write_o -> rmap_mem_nfee_comm_1:fee_0_rmap_write_i
	signal comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_rd_address_signal              : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_A:fee_codec_rmap_rd_address_o -> rmap_mem_nfee_comm_1:fee_0_rmap_rd_address_i
	signal rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_readdata_signal                      : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_1:fee_0_rmap_readdata_o -> COMM_Pedreiro_v1_01_A:fee_codec_rmap_readdata_i
	signal comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_wr_address_signal              : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_A:fee_codec_rmap_wr_address_o -> rmap_mem_nfee_comm_1:fee_0_rmap_wr_address_i
	signal comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_read_signal                    : std_logic;                      -- COMM_Pedreiro_v1_01_A:fee_codec_rmap_read_o -> rmap_mem_nfee_comm_1:fee_0_rmap_read_i
	signal rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_1:fee_0_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_A:fee_codec_rmap_wr_waitrequest_i
	signal comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_writedata_signal               : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_A:fee_codec_rmap_writedata_o -> rmap_mem_nfee_comm_1:fee_0_rmap_writedata_i
	signal rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_1:fee_0_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_A:fee_codec_rmap_rd_waitrequest_i
	signal comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_write_signal                   : std_logic;                      -- COMM_Pedreiro_v1_01_B:fee_codec_rmap_write_o -> rmap_mem_nfee_comm_2:fee_0_rmap_write_i
	signal comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_rd_address_signal              : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_B:fee_codec_rmap_rd_address_o -> rmap_mem_nfee_comm_2:fee_0_rmap_rd_address_i
	signal rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_readdata_signal                      : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_2:fee_0_rmap_readdata_o -> COMM_Pedreiro_v1_01_B:fee_codec_rmap_readdata_i
	signal comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_wr_address_signal              : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_B:fee_codec_rmap_wr_address_o -> rmap_mem_nfee_comm_2:fee_0_rmap_wr_address_i
	signal comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_read_signal                    : std_logic;                      -- COMM_Pedreiro_v1_01_B:fee_codec_rmap_read_o -> rmap_mem_nfee_comm_2:fee_0_rmap_read_i
	signal rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_2:fee_0_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_B:fee_codec_rmap_wr_waitrequest_i
	signal comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_writedata_signal               : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_B:fee_codec_rmap_writedata_o -> rmap_mem_nfee_comm_2:fee_0_rmap_writedata_i
	signal rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_2:fee_0_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_B:fee_codec_rmap_rd_waitrequest_i
	signal comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_write_signal                   : std_logic;                      -- COMM_Pedreiro_v1_01_D:fee_codec_rmap_write_o -> rmap_mem_nfee_comm_4:fee_0_rmap_write_i
	signal comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_rd_address_signal              : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_D:fee_codec_rmap_rd_address_o -> rmap_mem_nfee_comm_4:fee_0_rmap_rd_address_i
	signal rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_readdata_signal                      : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_4:fee_0_rmap_readdata_o -> COMM_Pedreiro_v1_01_D:fee_codec_rmap_readdata_i
	signal comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_wr_address_signal              : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_D:fee_codec_rmap_wr_address_o -> rmap_mem_nfee_comm_4:fee_0_rmap_wr_address_i
	signal comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_read_signal                    : std_logic;                      -- COMM_Pedreiro_v1_01_D:fee_codec_rmap_read_o -> rmap_mem_nfee_comm_4:fee_0_rmap_read_i
	signal rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_4:fee_0_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_D:fee_codec_rmap_wr_waitrequest_i
	signal comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_writedata_signal               : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_D:fee_codec_rmap_writedata_o -> rmap_mem_nfee_comm_4:fee_0_rmap_writedata_i
	signal rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_4:fee_0_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_D:fee_codec_rmap_rd_waitrequest_i
	signal comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_write_signal                   : std_logic;                      -- COMM_Pedreiro_v1_01_E:fee_codec_rmap_write_o -> rmap_mem_nfee_comm_5:fee_0_rmap_write_i
	signal comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_rd_address_signal              : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_E:fee_codec_rmap_rd_address_o -> rmap_mem_nfee_comm_5:fee_0_rmap_rd_address_i
	signal rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_readdata_signal                      : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_5:fee_0_rmap_readdata_o -> COMM_Pedreiro_v1_01_E:fee_codec_rmap_readdata_i
	signal comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_wr_address_signal              : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_E:fee_codec_rmap_wr_address_o -> rmap_mem_nfee_comm_5:fee_0_rmap_wr_address_i
	signal comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_read_signal                    : std_logic;                      -- COMM_Pedreiro_v1_01_E:fee_codec_rmap_read_o -> rmap_mem_nfee_comm_5:fee_0_rmap_read_i
	signal rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_5:fee_0_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_E:fee_codec_rmap_wr_waitrequest_i
	signal comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_writedata_signal               : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_E:fee_codec_rmap_writedata_o -> rmap_mem_nfee_comm_5:fee_0_rmap_writedata_i
	signal rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_5:fee_0_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_E:fee_codec_rmap_rd_waitrequest_i
	signal comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_write_signal                   : std_logic;                      -- COMM_Pedreiro_v1_01_F:fee_codec_rmap_write_o -> rmap_mem_nfee_comm_6:fee_0_rmap_write_i
	signal comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_rd_address_signal              : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_F:fee_codec_rmap_rd_address_o -> rmap_mem_nfee_comm_6:fee_0_rmap_rd_address_i
	signal rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_readdata_signal                      : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_6:fee_0_rmap_readdata_o -> COMM_Pedreiro_v1_01_F:fee_codec_rmap_readdata_i
	signal comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_wr_address_signal              : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_F:fee_codec_rmap_wr_address_o -> rmap_mem_nfee_comm_6:fee_0_rmap_wr_address_i
	signal comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_read_signal                    : std_logic;                      -- COMM_Pedreiro_v1_01_F:fee_codec_rmap_read_o -> rmap_mem_nfee_comm_6:fee_0_rmap_read_i
	signal rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_6:fee_0_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_F:fee_codec_rmap_wr_waitrequest_i
	signal comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_writedata_signal               : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_F:fee_codec_rmap_writedata_o -> rmap_mem_nfee_comm_6:fee_0_rmap_writedata_i
	signal rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_6:fee_0_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_F:fee_codec_rmap_rd_waitrequest_i
	signal comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_write_signal                      : std_logic;                      -- COMM_Pedreiro_v1_01_A:fee_hk_rmap_write_o -> rmap_mem_nfee_comm_1:fee_1_rmap_write_i
	signal comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_rd_address_signal                 : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_A:fee_hk_rmap_rd_address_o -> rmap_mem_nfee_comm_1:fee_1_rmap_rd_address_i
	signal rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_readdata_signal                      : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_1:fee_1_rmap_readdata_o -> COMM_Pedreiro_v1_01_A:fee_hk_rmap_readdata_i
	signal comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_wr_address_signal                 : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_A:fee_hk_rmap_wr_address_o -> rmap_mem_nfee_comm_1:fee_1_rmap_wr_address_i
	signal comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_read_signal                       : std_logic;                      -- COMM_Pedreiro_v1_01_A:fee_hk_rmap_read_o -> rmap_mem_nfee_comm_1:fee_1_rmap_read_i
	signal rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_1:fee_1_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_A:fee_hk_rmap_wr_waitrequest_i
	signal comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_writedata_signal                  : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_A:fee_hk_rmap_writedata_o -> rmap_mem_nfee_comm_1:fee_1_rmap_writedata_i
	signal rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_1:fee_1_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_A:fee_hk_rmap_rd_waitrequest_i
	signal comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_write_signal                      : std_logic;                      -- COMM_Pedreiro_v1_01_B:fee_hk_rmap_write_o -> rmap_mem_nfee_comm_2:fee_1_rmap_write_i
	signal comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_rd_address_signal                 : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_B:fee_hk_rmap_rd_address_o -> rmap_mem_nfee_comm_2:fee_1_rmap_rd_address_i
	signal rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_readdata_signal                      : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_2:fee_1_rmap_readdata_o -> COMM_Pedreiro_v1_01_B:fee_hk_rmap_readdata_i
	signal comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_wr_address_signal                 : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_B:fee_hk_rmap_wr_address_o -> rmap_mem_nfee_comm_2:fee_1_rmap_wr_address_i
	signal comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_read_signal                       : std_logic;                      -- COMM_Pedreiro_v1_01_B:fee_hk_rmap_read_o -> rmap_mem_nfee_comm_2:fee_1_rmap_read_i
	signal rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_2:fee_1_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_B:fee_hk_rmap_wr_waitrequest_i
	signal comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_writedata_signal                  : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_B:fee_hk_rmap_writedata_o -> rmap_mem_nfee_comm_2:fee_1_rmap_writedata_i
	signal rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_2:fee_1_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_B:fee_hk_rmap_rd_waitrequest_i
	signal comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_write_signal                      : std_logic;                      -- COMM_Pedreiro_v1_01_C:fee_hk_rmap_write_o -> rmap_mem_nfee_comm_3:fee_1_rmap_write_i
	signal comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_rd_address_signal                 : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_C:fee_hk_rmap_rd_address_o -> rmap_mem_nfee_comm_3:fee_1_rmap_rd_address_i
	signal rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_readdata_signal                      : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_3:fee_1_rmap_readdata_o -> COMM_Pedreiro_v1_01_C:fee_hk_rmap_readdata_i
	signal comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_wr_address_signal                 : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_C:fee_hk_rmap_wr_address_o -> rmap_mem_nfee_comm_3:fee_1_rmap_wr_address_i
	signal comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_read_signal                       : std_logic;                      -- COMM_Pedreiro_v1_01_C:fee_hk_rmap_read_o -> rmap_mem_nfee_comm_3:fee_1_rmap_read_i
	signal rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_3:fee_1_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_C:fee_hk_rmap_wr_waitrequest_i
	signal comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_writedata_signal                  : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_C:fee_hk_rmap_writedata_o -> rmap_mem_nfee_comm_3:fee_1_rmap_writedata_i
	signal rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_3:fee_1_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_C:fee_hk_rmap_rd_waitrequest_i
	signal comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_write_signal                      : std_logic;                      -- COMM_Pedreiro_v1_01_D:fee_hk_rmap_write_o -> rmap_mem_nfee_comm_4:fee_1_rmap_write_i
	signal comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_rd_address_signal                 : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_D:fee_hk_rmap_rd_address_o -> rmap_mem_nfee_comm_4:fee_1_rmap_rd_address_i
	signal rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_readdata_signal                      : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_4:fee_1_rmap_readdata_o -> COMM_Pedreiro_v1_01_D:fee_hk_rmap_readdata_i
	signal comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_wr_address_signal                 : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_D:fee_hk_rmap_wr_address_o -> rmap_mem_nfee_comm_4:fee_1_rmap_wr_address_i
	signal comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_read_signal                       : std_logic;                      -- COMM_Pedreiro_v1_01_D:fee_hk_rmap_read_o -> rmap_mem_nfee_comm_4:fee_1_rmap_read_i
	signal rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_4:fee_1_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_D:fee_hk_rmap_wr_waitrequest_i
	signal comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_writedata_signal                  : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_D:fee_hk_rmap_writedata_o -> rmap_mem_nfee_comm_4:fee_1_rmap_writedata_i
	signal rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_4:fee_1_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_D:fee_hk_rmap_rd_waitrequest_i
	signal comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_write_signal                      : std_logic;                      -- COMM_Pedreiro_v1_01_E:fee_hk_rmap_write_o -> rmap_mem_nfee_comm_5:fee_1_rmap_write_i
	signal comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_rd_address_signal                 : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_E:fee_hk_rmap_rd_address_o -> rmap_mem_nfee_comm_5:fee_1_rmap_rd_address_i
	signal rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_readdata_signal                      : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_5:fee_1_rmap_readdata_o -> COMM_Pedreiro_v1_01_E:fee_hk_rmap_readdata_i
	signal comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_wr_address_signal                 : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_E:fee_hk_rmap_wr_address_o -> rmap_mem_nfee_comm_5:fee_1_rmap_wr_address_i
	signal comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_read_signal                       : std_logic;                      -- COMM_Pedreiro_v1_01_E:fee_hk_rmap_read_o -> rmap_mem_nfee_comm_5:fee_1_rmap_read_i
	signal rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_5:fee_1_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_E:fee_hk_rmap_wr_waitrequest_i
	signal comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_writedata_signal                  : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_E:fee_hk_rmap_writedata_o -> rmap_mem_nfee_comm_5:fee_1_rmap_writedata_i
	signal rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_5:fee_1_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_E:fee_hk_rmap_rd_waitrequest_i
	signal comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_write_signal                      : std_logic;                      -- COMM_Pedreiro_v1_01_F:fee_hk_rmap_write_o -> rmap_mem_nfee_comm_6:fee_1_rmap_write_i
	signal comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_rd_address_signal                 : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_F:fee_hk_rmap_rd_address_o -> rmap_mem_nfee_comm_6:fee_1_rmap_rd_address_i
	signal rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_readdata_signal                      : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_6:fee_1_rmap_readdata_o -> COMM_Pedreiro_v1_01_F:fee_hk_rmap_readdata_i
	signal comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_wr_address_signal                 : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_F:fee_hk_rmap_wr_address_o -> rmap_mem_nfee_comm_6:fee_1_rmap_wr_address_i
	signal comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_read_signal                       : std_logic;                      -- COMM_Pedreiro_v1_01_F:fee_hk_rmap_read_o -> rmap_mem_nfee_comm_6:fee_1_rmap_read_i
	signal rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_6:fee_1_rmap_wr_waitrequest_o -> COMM_Pedreiro_v1_01_F:fee_hk_rmap_wr_waitrequest_i
	signal comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_writedata_signal                  : std_logic_vector(7 downto 0);   -- COMM_Pedreiro_v1_01_F:fee_hk_rmap_writedata_o -> rmap_mem_nfee_comm_6:fee_1_rmap_writedata_i
	signal rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal                : std_logic;                      -- rmap_mem_nfee_comm_6:fee_1_rmap_rd_waitrequest_o -> COMM_Pedreiro_v1_01_F:fee_hk_rmap_rd_waitrequest_i
	signal ext_flash_tcm_data_outen                                                               : std_logic;                      -- ext_flash:tcm_data_outen -> tristate_conduit_bridge_0:tcs_tcm_data_outen
	signal ext_flash_tcm_request                                                                  : std_logic;                      -- ext_flash:tcm_request -> tristate_conduit_bridge_0:request
	signal ext_flash_tcm_write_n_out                                                              : std_logic;                      -- ext_flash:tcm_write_n_out -> tristate_conduit_bridge_0:tcs_tcm_write_n_out
	signal ext_flash_tcm_read_n_out                                                               : std_logic;                      -- ext_flash:tcm_read_n_out -> tristate_conduit_bridge_0:tcs_tcm_read_n_out
	signal ext_flash_tcm_grant                                                                    : std_logic;                      -- tristate_conduit_bridge_0:grant -> ext_flash:tcm_grant
	signal ext_flash_tcm_chipselect_n_out                                                         : std_logic;                      -- ext_flash:tcm_chipselect_n_out -> tristate_conduit_bridge_0:tcs_tcm_chipselect_n_out
	signal ext_flash_tcm_address_out                                                              : std_logic_vector(25 downto 0);  -- ext_flash:tcm_address_out -> tristate_conduit_bridge_0:tcs_tcm_address_out
	signal ext_flash_tcm_data_out                                                                 : std_logic_vector(15 downto 0);  -- ext_flash:tcm_data_out -> tristate_conduit_bridge_0:tcs_tcm_data_out
	signal ext_flash_tcm_data_in                                                                  : std_logic_vector(15 downto 0);  -- tristate_conduit_bridge_0:tcs_tcm_data_in -> ext_flash:tcm_data_in
	signal rmap_mem_nfee_comm_1_avalon_mm_rmap_master_readdata                                    : std_logic_vector(7 downto 0);   -- mm_interconnect_0:rmap_mem_nfee_comm_1_avalon_mm_rmap_master_readdata -> rmap_mem_nfee_comm_1:avm_rmap_readdata_i
	signal rmap_mem_nfee_comm_1_avalon_mm_rmap_master_waitrequest                                 : std_logic;                      -- mm_interconnect_0:rmap_mem_nfee_comm_1_avalon_mm_rmap_master_waitrequest -> rmap_mem_nfee_comm_1:avm_rmap_waitrequest_i
	signal rmap_mem_nfee_comm_1_avalon_mm_rmap_master_address                                     : std_logic_vector(63 downto 0);  -- rmap_mem_nfee_comm_1:avm_rmap_address_o -> mm_interconnect_0:rmap_mem_nfee_comm_1_avalon_mm_rmap_master_address
	signal rmap_mem_nfee_comm_1_avalon_mm_rmap_master_read                                        : std_logic;                      -- rmap_mem_nfee_comm_1:avm_rmap_read_o -> mm_interconnect_0:rmap_mem_nfee_comm_1_avalon_mm_rmap_master_read
	signal rmap_mem_nfee_comm_1_avalon_mm_rmap_master_write                                       : std_logic;                      -- rmap_mem_nfee_comm_1:avm_rmap_write_o -> mm_interconnect_0:rmap_mem_nfee_comm_1_avalon_mm_rmap_master_write
	signal rmap_mem_nfee_comm_1_avalon_mm_rmap_master_writedata                                   : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_1:avm_rmap_writedata_o -> mm_interconnect_0:rmap_mem_nfee_comm_1_avalon_mm_rmap_master_writedata
	signal rmap_mem_nfee_comm_2_avalon_mm_rmap_master_readdata                                    : std_logic_vector(7 downto 0);   -- mm_interconnect_0:rmap_mem_nfee_comm_2_avalon_mm_rmap_master_readdata -> rmap_mem_nfee_comm_2:avm_rmap_readdata_i
	signal rmap_mem_nfee_comm_2_avalon_mm_rmap_master_waitrequest                                 : std_logic;                      -- mm_interconnect_0:rmap_mem_nfee_comm_2_avalon_mm_rmap_master_waitrequest -> rmap_mem_nfee_comm_2:avm_rmap_waitrequest_i
	signal rmap_mem_nfee_comm_2_avalon_mm_rmap_master_address                                     : std_logic_vector(63 downto 0);  -- rmap_mem_nfee_comm_2:avm_rmap_address_o -> mm_interconnect_0:rmap_mem_nfee_comm_2_avalon_mm_rmap_master_address
	signal rmap_mem_nfee_comm_2_avalon_mm_rmap_master_read                                        : std_logic;                      -- rmap_mem_nfee_comm_2:avm_rmap_read_o -> mm_interconnect_0:rmap_mem_nfee_comm_2_avalon_mm_rmap_master_read
	signal rmap_mem_nfee_comm_2_avalon_mm_rmap_master_write                                       : std_logic;                      -- rmap_mem_nfee_comm_2:avm_rmap_write_o -> mm_interconnect_0:rmap_mem_nfee_comm_2_avalon_mm_rmap_master_write
	signal rmap_mem_nfee_comm_2_avalon_mm_rmap_master_writedata                                   : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_2:avm_rmap_writedata_o -> mm_interconnect_0:rmap_mem_nfee_comm_2_avalon_mm_rmap_master_writedata
	signal rmap_mem_nfee_comm_3_avalon_mm_rmap_master_readdata                                    : std_logic_vector(7 downto 0);   -- mm_interconnect_0:rmap_mem_nfee_comm_3_avalon_mm_rmap_master_readdata -> rmap_mem_nfee_comm_3:avm_rmap_readdata_i
	signal rmap_mem_nfee_comm_3_avalon_mm_rmap_master_waitrequest                                 : std_logic;                      -- mm_interconnect_0:rmap_mem_nfee_comm_3_avalon_mm_rmap_master_waitrequest -> rmap_mem_nfee_comm_3:avm_rmap_waitrequest_i
	signal rmap_mem_nfee_comm_3_avalon_mm_rmap_master_address                                     : std_logic_vector(63 downto 0);  -- rmap_mem_nfee_comm_3:avm_rmap_address_o -> mm_interconnect_0:rmap_mem_nfee_comm_3_avalon_mm_rmap_master_address
	signal rmap_mem_nfee_comm_3_avalon_mm_rmap_master_read                                        : std_logic;                      -- rmap_mem_nfee_comm_3:avm_rmap_read_o -> mm_interconnect_0:rmap_mem_nfee_comm_3_avalon_mm_rmap_master_read
	signal rmap_mem_nfee_comm_3_avalon_mm_rmap_master_write                                       : std_logic;                      -- rmap_mem_nfee_comm_3:avm_rmap_write_o -> mm_interconnect_0:rmap_mem_nfee_comm_3_avalon_mm_rmap_master_write
	signal rmap_mem_nfee_comm_3_avalon_mm_rmap_master_writedata                                   : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_3:avm_rmap_writedata_o -> mm_interconnect_0:rmap_mem_nfee_comm_3_avalon_mm_rmap_master_writedata
	signal rmap_mem_nfee_comm_4_avalon_mm_rmap_master_readdata                                    : std_logic_vector(7 downto 0);   -- mm_interconnect_0:rmap_mem_nfee_comm_4_avalon_mm_rmap_master_readdata -> rmap_mem_nfee_comm_4:avm_rmap_readdata_i
	signal rmap_mem_nfee_comm_4_avalon_mm_rmap_master_waitrequest                                 : std_logic;                      -- mm_interconnect_0:rmap_mem_nfee_comm_4_avalon_mm_rmap_master_waitrequest -> rmap_mem_nfee_comm_4:avm_rmap_waitrequest_i
	signal rmap_mem_nfee_comm_4_avalon_mm_rmap_master_address                                     : std_logic_vector(63 downto 0);  -- rmap_mem_nfee_comm_4:avm_rmap_address_o -> mm_interconnect_0:rmap_mem_nfee_comm_4_avalon_mm_rmap_master_address
	signal rmap_mem_nfee_comm_4_avalon_mm_rmap_master_read                                        : std_logic;                      -- rmap_mem_nfee_comm_4:avm_rmap_read_o -> mm_interconnect_0:rmap_mem_nfee_comm_4_avalon_mm_rmap_master_read
	signal rmap_mem_nfee_comm_4_avalon_mm_rmap_master_write                                       : std_logic;                      -- rmap_mem_nfee_comm_4:avm_rmap_write_o -> mm_interconnect_0:rmap_mem_nfee_comm_4_avalon_mm_rmap_master_write
	signal rmap_mem_nfee_comm_4_avalon_mm_rmap_master_writedata                                   : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_4:avm_rmap_writedata_o -> mm_interconnect_0:rmap_mem_nfee_comm_4_avalon_mm_rmap_master_writedata
	signal rmap_mem_nfee_comm_5_avalon_mm_rmap_master_readdata                                    : std_logic_vector(7 downto 0);   -- mm_interconnect_0:rmap_mem_nfee_comm_5_avalon_mm_rmap_master_readdata -> rmap_mem_nfee_comm_5:avm_rmap_readdata_i
	signal rmap_mem_nfee_comm_5_avalon_mm_rmap_master_waitrequest                                 : std_logic;                      -- mm_interconnect_0:rmap_mem_nfee_comm_5_avalon_mm_rmap_master_waitrequest -> rmap_mem_nfee_comm_5:avm_rmap_waitrequest_i
	signal rmap_mem_nfee_comm_5_avalon_mm_rmap_master_address                                     : std_logic_vector(63 downto 0);  -- rmap_mem_nfee_comm_5:avm_rmap_address_o -> mm_interconnect_0:rmap_mem_nfee_comm_5_avalon_mm_rmap_master_address
	signal rmap_mem_nfee_comm_5_avalon_mm_rmap_master_read                                        : std_logic;                      -- rmap_mem_nfee_comm_5:avm_rmap_read_o -> mm_interconnect_0:rmap_mem_nfee_comm_5_avalon_mm_rmap_master_read
	signal rmap_mem_nfee_comm_5_avalon_mm_rmap_master_write                                       : std_logic;                      -- rmap_mem_nfee_comm_5:avm_rmap_write_o -> mm_interconnect_0:rmap_mem_nfee_comm_5_avalon_mm_rmap_master_write
	signal rmap_mem_nfee_comm_5_avalon_mm_rmap_master_writedata                                   : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_5:avm_rmap_writedata_o -> mm_interconnect_0:rmap_mem_nfee_comm_5_avalon_mm_rmap_master_writedata
	signal rmap_mem_nfee_comm_6_avalon_mm_rmap_master_readdata                                    : std_logic_vector(7 downto 0);   -- mm_interconnect_0:rmap_mem_nfee_comm_6_avalon_mm_rmap_master_readdata -> rmap_mem_nfee_comm_6:avm_rmap_readdata_i
	signal rmap_mem_nfee_comm_6_avalon_mm_rmap_master_waitrequest                                 : std_logic;                      -- mm_interconnect_0:rmap_mem_nfee_comm_6_avalon_mm_rmap_master_waitrequest -> rmap_mem_nfee_comm_6:avm_rmap_waitrequest_i
	signal rmap_mem_nfee_comm_6_avalon_mm_rmap_master_address                                     : std_logic_vector(63 downto 0);  -- rmap_mem_nfee_comm_6:avm_rmap_address_o -> mm_interconnect_0:rmap_mem_nfee_comm_6_avalon_mm_rmap_master_address
	signal rmap_mem_nfee_comm_6_avalon_mm_rmap_master_read                                        : std_logic;                      -- rmap_mem_nfee_comm_6:avm_rmap_read_o -> mm_interconnect_0:rmap_mem_nfee_comm_6_avalon_mm_rmap_master_read
	signal rmap_mem_nfee_comm_6_avalon_mm_rmap_master_write                                       : std_logic;                      -- rmap_mem_nfee_comm_6:avm_rmap_write_o -> mm_interconnect_0:rmap_mem_nfee_comm_6_avalon_mm_rmap_master_write
	signal rmap_mem_nfee_comm_6_avalon_mm_rmap_master_writedata                                   : std_logic_vector(7 downto 0);   -- rmap_mem_nfee_comm_6:avm_rmap_writedata_o -> mm_interconnect_0:rmap_mem_nfee_comm_6_avalon_mm_rmap_master_writedata
	signal ddr2_address_span_extender_expanded_master_waitrequest                                 : std_logic;                      -- mm_interconnect_0:ddr2_address_span_extender_expanded_master_waitrequest -> ddr2_address_span_extender:avm_m0_waitrequest
	signal ddr2_address_span_extender_expanded_master_readdata                                    : std_logic_vector(31 downto 0);  -- mm_interconnect_0:ddr2_address_span_extender_expanded_master_readdata -> ddr2_address_span_extender:avm_m0_readdata
	signal ddr2_address_span_extender_expanded_master_address                                     : std_logic_vector(31 downto 0);  -- ddr2_address_span_extender:avm_m0_address -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_address
	signal ddr2_address_span_extender_expanded_master_read                                        : std_logic;                      -- ddr2_address_span_extender:avm_m0_read -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_read
	signal ddr2_address_span_extender_expanded_master_byteenable                                  : std_logic_vector(3 downto 0);   -- ddr2_address_span_extender:avm_m0_byteenable -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_byteenable
	signal ddr2_address_span_extender_expanded_master_readdatavalid                               : std_logic;                      -- mm_interconnect_0:ddr2_address_span_extender_expanded_master_readdatavalid -> ddr2_address_span_extender:avm_m0_readdatavalid
	signal ddr2_address_span_extender_expanded_master_write                                       : std_logic;                      -- ddr2_address_span_extender:avm_m0_write -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_write
	signal ddr2_address_span_extender_expanded_master_writedata                                   : std_logic_vector(31 downto 0);  -- ddr2_address_span_extender:avm_m0_writedata -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_writedata
	signal ddr2_address_span_extender_expanded_master_burstcount                                  : std_logic_vector(7 downto 0);   -- ddr2_address_span_extender:avm_m0_burstcount -> mm_interconnect_0:ddr2_address_span_extender_expanded_master_burstcount
	signal dma_comm_1_left_mm_read_readdata                                                       : std_logic_vector(255 downto 0); -- mm_interconnect_0:dma_comm_1_left_mm_read_readdata -> dma_comm_1_left:mm_read_readdata
	signal dma_comm_1_left_mm_read_waitrequest                                                    : std_logic;                      -- mm_interconnect_0:dma_comm_1_left_mm_read_waitrequest -> dma_comm_1_left:mm_read_waitrequest
	signal dma_comm_1_left_mm_read_address                                                        : std_logic_vector(31 downto 0);  -- dma_comm_1_left:mm_read_address -> mm_interconnect_0:dma_comm_1_left_mm_read_address
	signal dma_comm_1_left_mm_read_read                                                           : std_logic;                      -- dma_comm_1_left:mm_read_read -> mm_interconnect_0:dma_comm_1_left_mm_read_read
	signal dma_comm_1_left_mm_read_byteenable                                                     : std_logic_vector(31 downto 0);  -- dma_comm_1_left:mm_read_byteenable -> mm_interconnect_0:dma_comm_1_left_mm_read_byteenable
	signal dma_comm_1_left_mm_read_readdatavalid                                                  : std_logic;                      -- mm_interconnect_0:dma_comm_1_left_mm_read_readdatavalid -> dma_comm_1_left:mm_read_readdatavalid
	signal dma_comm_6_right_mm_read_readdata                                                      : std_logic_vector(255 downto 0); -- mm_interconnect_0:dma_comm_6_right_mm_read_readdata -> dma_comm_6_right:mm_read_readdata
	signal dma_comm_6_right_mm_read_waitrequest                                                   : std_logic;                      -- mm_interconnect_0:dma_comm_6_right_mm_read_waitrequest -> dma_comm_6_right:mm_read_waitrequest
	signal dma_comm_6_right_mm_read_address                                                       : std_logic_vector(31 downto 0);  -- dma_comm_6_right:mm_read_address -> mm_interconnect_0:dma_comm_6_right_mm_read_address
	signal dma_comm_6_right_mm_read_read                                                          : std_logic;                      -- dma_comm_6_right:mm_read_read -> mm_interconnect_0:dma_comm_6_right_mm_read_read
	signal dma_comm_6_right_mm_read_byteenable                                                    : std_logic_vector(31 downto 0);  -- dma_comm_6_right:mm_read_byteenable -> mm_interconnect_0:dma_comm_6_right_mm_read_byteenable
	signal dma_comm_6_right_mm_read_readdatavalid                                                 : std_logic;                      -- mm_interconnect_0:dma_comm_6_right_mm_read_readdatavalid -> dma_comm_6_right:mm_read_readdatavalid
	signal dma_comm_6_left_mm_read_readdata                                                       : std_logic_vector(255 downto 0); -- mm_interconnect_0:dma_comm_6_left_mm_read_readdata -> dma_comm_6_left:mm_read_readdata
	signal dma_comm_6_left_mm_read_waitrequest                                                    : std_logic;                      -- mm_interconnect_0:dma_comm_6_left_mm_read_waitrequest -> dma_comm_6_left:mm_read_waitrequest
	signal dma_comm_6_left_mm_read_address                                                        : std_logic_vector(31 downto 0);  -- dma_comm_6_left:mm_read_address -> mm_interconnect_0:dma_comm_6_left_mm_read_address
	signal dma_comm_6_left_mm_read_read                                                           : std_logic;                      -- dma_comm_6_left:mm_read_read -> mm_interconnect_0:dma_comm_6_left_mm_read_read
	signal dma_comm_6_left_mm_read_byteenable                                                     : std_logic_vector(31 downto 0);  -- dma_comm_6_left:mm_read_byteenable -> mm_interconnect_0:dma_comm_6_left_mm_read_byteenable
	signal dma_comm_6_left_mm_read_readdatavalid                                                  : std_logic;                      -- mm_interconnect_0:dma_comm_6_left_mm_read_readdatavalid -> dma_comm_6_left:mm_read_readdatavalid
	signal dma_comm_5_right_mm_read_readdata                                                      : std_logic_vector(255 downto 0); -- mm_interconnect_0:dma_comm_5_right_mm_read_readdata -> dma_comm_5_right:mm_read_readdata
	signal dma_comm_5_right_mm_read_waitrequest                                                   : std_logic;                      -- mm_interconnect_0:dma_comm_5_right_mm_read_waitrequest -> dma_comm_5_right:mm_read_waitrequest
	signal dma_comm_5_right_mm_read_address                                                       : std_logic_vector(31 downto 0);  -- dma_comm_5_right:mm_read_address -> mm_interconnect_0:dma_comm_5_right_mm_read_address
	signal dma_comm_5_right_mm_read_read                                                          : std_logic;                      -- dma_comm_5_right:mm_read_read -> mm_interconnect_0:dma_comm_5_right_mm_read_read
	signal dma_comm_5_right_mm_read_byteenable                                                    : std_logic_vector(31 downto 0);  -- dma_comm_5_right:mm_read_byteenable -> mm_interconnect_0:dma_comm_5_right_mm_read_byteenable
	signal dma_comm_5_right_mm_read_readdatavalid                                                 : std_logic;                      -- mm_interconnect_0:dma_comm_5_right_mm_read_readdatavalid -> dma_comm_5_right:mm_read_readdatavalid
	signal dma_comm_5_left_mm_read_readdata                                                       : std_logic_vector(255 downto 0); -- mm_interconnect_0:dma_comm_5_left_mm_read_readdata -> dma_comm_5_left:mm_read_readdata
	signal dma_comm_5_left_mm_read_waitrequest                                                    : std_logic;                      -- mm_interconnect_0:dma_comm_5_left_mm_read_waitrequest -> dma_comm_5_left:mm_read_waitrequest
	signal dma_comm_5_left_mm_read_address                                                        : std_logic_vector(31 downto 0);  -- dma_comm_5_left:mm_read_address -> mm_interconnect_0:dma_comm_5_left_mm_read_address
	signal dma_comm_5_left_mm_read_read                                                           : std_logic;                      -- dma_comm_5_left:mm_read_read -> mm_interconnect_0:dma_comm_5_left_mm_read_read
	signal dma_comm_5_left_mm_read_byteenable                                                     : std_logic_vector(31 downto 0);  -- dma_comm_5_left:mm_read_byteenable -> mm_interconnect_0:dma_comm_5_left_mm_read_byteenable
	signal dma_comm_5_left_mm_read_readdatavalid                                                  : std_logic;                      -- mm_interconnect_0:dma_comm_5_left_mm_read_readdatavalid -> dma_comm_5_left:mm_read_readdatavalid
	signal dma_comm_4_right_mm_read_readdata                                                      : std_logic_vector(255 downto 0); -- mm_interconnect_0:dma_comm_4_right_mm_read_readdata -> dma_comm_4_right:mm_read_readdata
	signal dma_comm_4_right_mm_read_waitrequest                                                   : std_logic;                      -- mm_interconnect_0:dma_comm_4_right_mm_read_waitrequest -> dma_comm_4_right:mm_read_waitrequest
	signal dma_comm_4_right_mm_read_address                                                       : std_logic_vector(31 downto 0);  -- dma_comm_4_right:mm_read_address -> mm_interconnect_0:dma_comm_4_right_mm_read_address
	signal dma_comm_4_right_mm_read_read                                                          : std_logic;                      -- dma_comm_4_right:mm_read_read -> mm_interconnect_0:dma_comm_4_right_mm_read_read
	signal dma_comm_4_right_mm_read_byteenable                                                    : std_logic_vector(31 downto 0);  -- dma_comm_4_right:mm_read_byteenable -> mm_interconnect_0:dma_comm_4_right_mm_read_byteenable
	signal dma_comm_4_right_mm_read_readdatavalid                                                 : std_logic;                      -- mm_interconnect_0:dma_comm_4_right_mm_read_readdatavalid -> dma_comm_4_right:mm_read_readdatavalid
	signal dma_comm_4_left_mm_read_readdata                                                       : std_logic_vector(255 downto 0); -- mm_interconnect_0:dma_comm_4_left_mm_read_readdata -> dma_comm_4_left:mm_read_readdata
	signal dma_comm_4_left_mm_read_waitrequest                                                    : std_logic;                      -- mm_interconnect_0:dma_comm_4_left_mm_read_waitrequest -> dma_comm_4_left:mm_read_waitrequest
	signal dma_comm_4_left_mm_read_address                                                        : std_logic_vector(31 downto 0);  -- dma_comm_4_left:mm_read_address -> mm_interconnect_0:dma_comm_4_left_mm_read_address
	signal dma_comm_4_left_mm_read_read                                                           : std_logic;                      -- dma_comm_4_left:mm_read_read -> mm_interconnect_0:dma_comm_4_left_mm_read_read
	signal dma_comm_4_left_mm_read_byteenable                                                     : std_logic_vector(31 downto 0);  -- dma_comm_4_left:mm_read_byteenable -> mm_interconnect_0:dma_comm_4_left_mm_read_byteenable
	signal dma_comm_4_left_mm_read_readdatavalid                                                  : std_logic;                      -- mm_interconnect_0:dma_comm_4_left_mm_read_readdatavalid -> dma_comm_4_left:mm_read_readdatavalid
	signal dma_comm_3_right_mm_read_readdata                                                      : std_logic_vector(255 downto 0); -- mm_interconnect_0:dma_comm_3_right_mm_read_readdata -> dma_comm_3_right:mm_read_readdata
	signal dma_comm_3_right_mm_read_waitrequest                                                   : std_logic;                      -- mm_interconnect_0:dma_comm_3_right_mm_read_waitrequest -> dma_comm_3_right:mm_read_waitrequest
	signal dma_comm_3_right_mm_read_address                                                       : std_logic_vector(31 downto 0);  -- dma_comm_3_right:mm_read_address -> mm_interconnect_0:dma_comm_3_right_mm_read_address
	signal dma_comm_3_right_mm_read_read                                                          : std_logic;                      -- dma_comm_3_right:mm_read_read -> mm_interconnect_0:dma_comm_3_right_mm_read_read
	signal dma_comm_3_right_mm_read_byteenable                                                    : std_logic_vector(31 downto 0);  -- dma_comm_3_right:mm_read_byteenable -> mm_interconnect_0:dma_comm_3_right_mm_read_byteenable
	signal dma_comm_3_right_mm_read_readdatavalid                                                 : std_logic;                      -- mm_interconnect_0:dma_comm_3_right_mm_read_readdatavalid -> dma_comm_3_right:mm_read_readdatavalid
	signal dma_comm_3_left_mm_read_readdata                                                       : std_logic_vector(255 downto 0); -- mm_interconnect_0:dma_comm_3_left_mm_read_readdata -> dma_comm_3_left:mm_read_readdata
	signal dma_comm_3_left_mm_read_waitrequest                                                    : std_logic;                      -- mm_interconnect_0:dma_comm_3_left_mm_read_waitrequest -> dma_comm_3_left:mm_read_waitrequest
	signal dma_comm_3_left_mm_read_address                                                        : std_logic_vector(31 downto 0);  -- dma_comm_3_left:mm_read_address -> mm_interconnect_0:dma_comm_3_left_mm_read_address
	signal dma_comm_3_left_mm_read_read                                                           : std_logic;                      -- dma_comm_3_left:mm_read_read -> mm_interconnect_0:dma_comm_3_left_mm_read_read
	signal dma_comm_3_left_mm_read_byteenable                                                     : std_logic_vector(31 downto 0);  -- dma_comm_3_left:mm_read_byteenable -> mm_interconnect_0:dma_comm_3_left_mm_read_byteenable
	signal dma_comm_3_left_mm_read_readdatavalid                                                  : std_logic;                      -- mm_interconnect_0:dma_comm_3_left_mm_read_readdatavalid -> dma_comm_3_left:mm_read_readdatavalid
	signal dma_comm_2_right_mm_read_readdata                                                      : std_logic_vector(255 downto 0); -- mm_interconnect_0:dma_comm_2_right_mm_read_readdata -> dma_comm_2_right:mm_read_readdata
	signal dma_comm_2_right_mm_read_waitrequest                                                   : std_logic;                      -- mm_interconnect_0:dma_comm_2_right_mm_read_waitrequest -> dma_comm_2_right:mm_read_waitrequest
	signal dma_comm_2_right_mm_read_address                                                       : std_logic_vector(31 downto 0);  -- dma_comm_2_right:mm_read_address -> mm_interconnect_0:dma_comm_2_right_mm_read_address
	signal dma_comm_2_right_mm_read_read                                                          : std_logic;                      -- dma_comm_2_right:mm_read_read -> mm_interconnect_0:dma_comm_2_right_mm_read_read
	signal dma_comm_2_right_mm_read_byteenable                                                    : std_logic_vector(31 downto 0);  -- dma_comm_2_right:mm_read_byteenable -> mm_interconnect_0:dma_comm_2_right_mm_read_byteenable
	signal dma_comm_2_right_mm_read_readdatavalid                                                 : std_logic;                      -- mm_interconnect_0:dma_comm_2_right_mm_read_readdatavalid -> dma_comm_2_right:mm_read_readdatavalid
	signal dma_comm_2_left_mm_read_readdata                                                       : std_logic_vector(255 downto 0); -- mm_interconnect_0:dma_comm_2_left_mm_read_readdata -> dma_comm_2_left:mm_read_readdata
	signal dma_comm_2_left_mm_read_waitrequest                                                    : std_logic;                      -- mm_interconnect_0:dma_comm_2_left_mm_read_waitrequest -> dma_comm_2_left:mm_read_waitrequest
	signal dma_comm_2_left_mm_read_address                                                        : std_logic_vector(31 downto 0);  -- dma_comm_2_left:mm_read_address -> mm_interconnect_0:dma_comm_2_left_mm_read_address
	signal dma_comm_2_left_mm_read_read                                                           : std_logic;                      -- dma_comm_2_left:mm_read_read -> mm_interconnect_0:dma_comm_2_left_mm_read_read
	signal dma_comm_2_left_mm_read_byteenable                                                     : std_logic_vector(31 downto 0);  -- dma_comm_2_left:mm_read_byteenable -> mm_interconnect_0:dma_comm_2_left_mm_read_byteenable
	signal dma_comm_2_left_mm_read_readdatavalid                                                  : std_logic;                      -- mm_interconnect_0:dma_comm_2_left_mm_read_readdatavalid -> dma_comm_2_left:mm_read_readdatavalid
	signal dma_comm_1_right_mm_read_readdata                                                      : std_logic_vector(255 downto 0); -- mm_interconnect_0:dma_comm_1_right_mm_read_readdata -> dma_comm_1_right:mm_read_readdata
	signal dma_comm_1_right_mm_read_waitrequest                                                   : std_logic;                      -- mm_interconnect_0:dma_comm_1_right_mm_read_waitrequest -> dma_comm_1_right:mm_read_waitrequest
	signal dma_comm_1_right_mm_read_address                                                       : std_logic_vector(31 downto 0);  -- dma_comm_1_right:mm_read_address -> mm_interconnect_0:dma_comm_1_right_mm_read_address
	signal dma_comm_1_right_mm_read_read                                                          : std_logic;                      -- dma_comm_1_right:mm_read_read -> mm_interconnect_0:dma_comm_1_right_mm_read_read
	signal dma_comm_1_right_mm_read_byteenable                                                    : std_logic_vector(31 downto 0);  -- dma_comm_1_right:mm_read_byteenable -> mm_interconnect_0:dma_comm_1_right_mm_read_byteenable
	signal dma_comm_1_right_mm_read_readdatavalid                                                 : std_logic;                      -- mm_interconnect_0:dma_comm_1_right_mm_read_readdatavalid -> dma_comm_1_right:mm_read_readdatavalid
	signal dma_ftdi_usb3_mm_write_waitrequest                                                     : std_logic;                      -- mm_interconnect_0:dma_ftdi_usb3_mm_write_waitrequest -> dma_ftdi_usb3:mm_write_waitrequest
	signal dma_ftdi_usb3_mm_write_address                                                         : std_logic_vector(31 downto 0);  -- dma_ftdi_usb3:mm_write_address -> mm_interconnect_0:dma_ftdi_usb3_mm_write_address
	signal dma_ftdi_usb3_mm_write_byteenable                                                      : std_logic_vector(31 downto 0);  -- dma_ftdi_usb3:mm_write_byteenable -> mm_interconnect_0:dma_ftdi_usb3_mm_write_byteenable
	signal dma_ftdi_usb3_mm_write_write                                                           : std_logic;                      -- dma_ftdi_usb3:mm_write_write -> mm_interconnect_0:dma_ftdi_usb3_mm_write_write
	signal dma_ftdi_usb3_mm_write_writedata                                                       : std_logic_vector(255 downto 0); -- dma_ftdi_usb3:mm_write_writedata -> mm_interconnect_0:dma_ftdi_usb3_mm_write_writedata
	signal mm_interconnect_0_m2_ddr2_memory_avl_beginbursttransfer                                : std_logic;                      -- mm_interconnect_0:m2_ddr2_memory_avl_beginbursttransfer -> m2_ddr2_memory:avl_burstbegin
	signal mm_interconnect_0_m2_ddr2_memory_avl_readdata                                          : std_logic_vector(255 downto 0); -- m2_ddr2_memory:avl_rdata -> mm_interconnect_0:m2_ddr2_memory_avl_readdata
	signal m2_ddr2_memory_avl_waitrequest                                                         : std_logic;                      -- m2_ddr2_memory:avl_ready -> m2_ddr2_memory_avl_waitrequest:in
	signal mm_interconnect_0_m2_ddr2_memory_avl_address                                           : std_logic_vector(25 downto 0);  -- mm_interconnect_0:m2_ddr2_memory_avl_address -> m2_ddr2_memory:avl_addr
	signal mm_interconnect_0_m2_ddr2_memory_avl_read                                              : std_logic;                      -- mm_interconnect_0:m2_ddr2_memory_avl_read -> m2_ddr2_memory:avl_read_req
	signal mm_interconnect_0_m2_ddr2_memory_avl_byteenable                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_0:m2_ddr2_memory_avl_byteenable -> m2_ddr2_memory:avl_be
	signal mm_interconnect_0_m2_ddr2_memory_avl_readdatavalid                                     : std_logic;                      -- m2_ddr2_memory:avl_rdata_valid -> mm_interconnect_0:m2_ddr2_memory_avl_readdatavalid
	signal mm_interconnect_0_m2_ddr2_memory_avl_write                                             : std_logic;                      -- mm_interconnect_0:m2_ddr2_memory_avl_write -> m2_ddr2_memory:avl_write_req
	signal mm_interconnect_0_m2_ddr2_memory_avl_writedata                                         : std_logic_vector(255 downto 0); -- mm_interconnect_0:m2_ddr2_memory_avl_writedata -> m2_ddr2_memory:avl_wdata
	signal mm_interconnect_0_m2_ddr2_memory_avl_burstcount                                        : std_logic_vector(7 downto 0);   -- mm_interconnect_0:m2_ddr2_memory_avl_burstcount -> m2_ddr2_memory:avl_size
	signal mm_interconnect_0_m1_clock_bridge_s0_readdata                                          : std_logic_vector(255 downto 0); -- m1_clock_bridge:s0_readdata -> mm_interconnect_0:m1_clock_bridge_s0_readdata
	signal mm_interconnect_0_m1_clock_bridge_s0_waitrequest                                       : std_logic;                      -- m1_clock_bridge:s0_waitrequest -> mm_interconnect_0:m1_clock_bridge_s0_waitrequest
	signal mm_interconnect_0_m1_clock_bridge_s0_debugaccess                                       : std_logic;                      -- mm_interconnect_0:m1_clock_bridge_s0_debugaccess -> m1_clock_bridge:s0_debugaccess
	signal mm_interconnect_0_m1_clock_bridge_s0_address                                           : std_logic_vector(30 downto 0);  -- mm_interconnect_0:m1_clock_bridge_s0_address -> m1_clock_bridge:s0_address
	signal mm_interconnect_0_m1_clock_bridge_s0_read                                              : std_logic;                      -- mm_interconnect_0:m1_clock_bridge_s0_read -> m1_clock_bridge:s0_read
	signal mm_interconnect_0_m1_clock_bridge_s0_byteenable                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_0:m1_clock_bridge_s0_byteenable -> m1_clock_bridge:s0_byteenable
	signal mm_interconnect_0_m1_clock_bridge_s0_readdatavalid                                     : std_logic;                      -- m1_clock_bridge:s0_readdatavalid -> mm_interconnect_0:m1_clock_bridge_s0_readdatavalid
	signal mm_interconnect_0_m1_clock_bridge_s0_write                                             : std_logic;                      -- mm_interconnect_0:m1_clock_bridge_s0_write -> m1_clock_bridge:s0_write
	signal mm_interconnect_0_m1_clock_bridge_s0_writedata                                         : std_logic_vector(255 downto 0); -- mm_interconnect_0:m1_clock_bridge_s0_writedata -> m1_clock_bridge:s0_writedata
	signal mm_interconnect_0_m1_clock_bridge_s0_burstcount                                        : std_logic_vector(2 downto 0);   -- mm_interconnect_0:m1_clock_bridge_s0_burstcount -> m1_clock_bridge:s0_burstcount
	signal nios2_gen2_0_data_master_readdata                                                      : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                                   : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                                   : std_logic;                      -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                                       : std_logic_vector(31 downto 0);  -- nios2_gen2_0:d_address -> mm_interconnect_1:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                                    : std_logic_vector(3 downto 0);   -- nios2_gen2_0:d_byteenable -> mm_interconnect_1:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                                          : std_logic;                      -- nios2_gen2_0:d_read -> mm_interconnect_1:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                                         : std_logic;                      -- nios2_gen2_0:d_write -> mm_interconnect_1:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                                     : std_logic_vector(31 downto 0);  -- nios2_gen2_0:d_writedata -> mm_interconnect_1:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                                               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                                            : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                                                : std_logic_vector(31 downto 0);  -- nios2_gen2_0:i_address -> mm_interconnect_1:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                                   : std_logic;                      -- nios2_gen2_0:i_read -> mm_interconnect_1:nios2_gen2_0_instruction_master_read
	signal nios2_gen2_0_instruction_master_readdatavalid                                          : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	signal nios2_gen2_0_instruction_master_burstcount                                             : std_logic_vector(3 downto 0);   -- nios2_gen2_0:i_burstcount -> mm_interconnect_1:nios2_gen2_0_instruction_master_burstcount
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect                             : std_logic;                      -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata                               : std_logic_vector(31 downto 0);  -- jtag_uart_0:av_readdata -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest                            : std_logic;                      -- jtag_uart_0:av_waitrequest -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address                                : std_logic_vector(0 downto 0);   -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read                                   : std_logic;                      -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write                                  : std_logic;                      -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata                              : std_logic_vector(31 downto 0);  -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_readdata                    : std_logic_vector(31 downto 0);  -- rmap_mem_nfee_comm_1:avs_0_rmap_readdata_o -> mm_interconnect_1:rmap_mem_nfee_comm_1_avalon_rmap_slave_0_readdata
	signal mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_waitrequest                 : std_logic;                      -- rmap_mem_nfee_comm_1:avs_0_rmap_waitrequest_o -> mm_interconnect_1:rmap_mem_nfee_comm_1_avalon_rmap_slave_0_waitrequest
	signal mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_address                     : std_logic_vector(11 downto 0);  -- mm_interconnect_1:rmap_mem_nfee_comm_1_avalon_rmap_slave_0_address -> rmap_mem_nfee_comm_1:avs_0_rmap_address_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_read                        : std_logic;                      -- mm_interconnect_1:rmap_mem_nfee_comm_1_avalon_rmap_slave_0_read -> rmap_mem_nfee_comm_1:avs_0_rmap_read_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_byteenable                  : std_logic_vector(3 downto 0);   -- mm_interconnect_1:rmap_mem_nfee_comm_1_avalon_rmap_slave_0_byteenable -> rmap_mem_nfee_comm_1:avs_0_rmap_byteenable_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_write                       : std_logic;                      -- mm_interconnect_1:rmap_mem_nfee_comm_1_avalon_rmap_slave_0_write -> rmap_mem_nfee_comm_1:avs_0_rmap_write_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:rmap_mem_nfee_comm_1_avalon_rmap_slave_0_writedata -> rmap_mem_nfee_comm_1:avs_0_rmap_writedata_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_readdata                    : std_logic_vector(31 downto 0);  -- rmap_mem_nfee_comm_2:avs_0_rmap_readdata_o -> mm_interconnect_1:rmap_mem_nfee_comm_2_avalon_rmap_slave_0_readdata
	signal mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_waitrequest                 : std_logic;                      -- rmap_mem_nfee_comm_2:avs_0_rmap_waitrequest_o -> mm_interconnect_1:rmap_mem_nfee_comm_2_avalon_rmap_slave_0_waitrequest
	signal mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_address                     : std_logic_vector(11 downto 0);  -- mm_interconnect_1:rmap_mem_nfee_comm_2_avalon_rmap_slave_0_address -> rmap_mem_nfee_comm_2:avs_0_rmap_address_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_read                        : std_logic;                      -- mm_interconnect_1:rmap_mem_nfee_comm_2_avalon_rmap_slave_0_read -> rmap_mem_nfee_comm_2:avs_0_rmap_read_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_byteenable                  : std_logic_vector(3 downto 0);   -- mm_interconnect_1:rmap_mem_nfee_comm_2_avalon_rmap_slave_0_byteenable -> rmap_mem_nfee_comm_2:avs_0_rmap_byteenable_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_write                       : std_logic;                      -- mm_interconnect_1:rmap_mem_nfee_comm_2_avalon_rmap_slave_0_write -> rmap_mem_nfee_comm_2:avs_0_rmap_write_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:rmap_mem_nfee_comm_2_avalon_rmap_slave_0_writedata -> rmap_mem_nfee_comm_2:avs_0_rmap_writedata_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_readdata                    : std_logic_vector(31 downto 0);  -- rmap_mem_nfee_comm_3:avs_0_rmap_readdata_o -> mm_interconnect_1:rmap_mem_nfee_comm_3_avalon_rmap_slave_0_readdata
	signal mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_waitrequest                 : std_logic;                      -- rmap_mem_nfee_comm_3:avs_0_rmap_waitrequest_o -> mm_interconnect_1:rmap_mem_nfee_comm_3_avalon_rmap_slave_0_waitrequest
	signal mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_address                     : std_logic_vector(11 downto 0);  -- mm_interconnect_1:rmap_mem_nfee_comm_3_avalon_rmap_slave_0_address -> rmap_mem_nfee_comm_3:avs_0_rmap_address_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_read                        : std_logic;                      -- mm_interconnect_1:rmap_mem_nfee_comm_3_avalon_rmap_slave_0_read -> rmap_mem_nfee_comm_3:avs_0_rmap_read_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_byteenable                  : std_logic_vector(3 downto 0);   -- mm_interconnect_1:rmap_mem_nfee_comm_3_avalon_rmap_slave_0_byteenable -> rmap_mem_nfee_comm_3:avs_0_rmap_byteenable_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_write                       : std_logic;                      -- mm_interconnect_1:rmap_mem_nfee_comm_3_avalon_rmap_slave_0_write -> rmap_mem_nfee_comm_3:avs_0_rmap_write_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:rmap_mem_nfee_comm_3_avalon_rmap_slave_0_writedata -> rmap_mem_nfee_comm_3:avs_0_rmap_writedata_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_readdata                    : std_logic_vector(31 downto 0);  -- rmap_mem_nfee_comm_4:avs_0_rmap_readdata_o -> mm_interconnect_1:rmap_mem_nfee_comm_4_avalon_rmap_slave_0_readdata
	signal mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_waitrequest                 : std_logic;                      -- rmap_mem_nfee_comm_4:avs_0_rmap_waitrequest_o -> mm_interconnect_1:rmap_mem_nfee_comm_4_avalon_rmap_slave_0_waitrequest
	signal mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_address                     : std_logic_vector(11 downto 0);  -- mm_interconnect_1:rmap_mem_nfee_comm_4_avalon_rmap_slave_0_address -> rmap_mem_nfee_comm_4:avs_0_rmap_address_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_read                        : std_logic;                      -- mm_interconnect_1:rmap_mem_nfee_comm_4_avalon_rmap_slave_0_read -> rmap_mem_nfee_comm_4:avs_0_rmap_read_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_byteenable                  : std_logic_vector(3 downto 0);   -- mm_interconnect_1:rmap_mem_nfee_comm_4_avalon_rmap_slave_0_byteenable -> rmap_mem_nfee_comm_4:avs_0_rmap_byteenable_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_write                       : std_logic;                      -- mm_interconnect_1:rmap_mem_nfee_comm_4_avalon_rmap_slave_0_write -> rmap_mem_nfee_comm_4:avs_0_rmap_write_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:rmap_mem_nfee_comm_4_avalon_rmap_slave_0_writedata -> rmap_mem_nfee_comm_4:avs_0_rmap_writedata_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_readdata                    : std_logic_vector(31 downto 0);  -- rmap_mem_nfee_comm_5:avs_0_rmap_readdata_o -> mm_interconnect_1:rmap_mem_nfee_comm_5_avalon_rmap_slave_0_readdata
	signal mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_waitrequest                 : std_logic;                      -- rmap_mem_nfee_comm_5:avs_0_rmap_waitrequest_o -> mm_interconnect_1:rmap_mem_nfee_comm_5_avalon_rmap_slave_0_waitrequest
	signal mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_address                     : std_logic_vector(11 downto 0);  -- mm_interconnect_1:rmap_mem_nfee_comm_5_avalon_rmap_slave_0_address -> rmap_mem_nfee_comm_5:avs_0_rmap_address_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_read                        : std_logic;                      -- mm_interconnect_1:rmap_mem_nfee_comm_5_avalon_rmap_slave_0_read -> rmap_mem_nfee_comm_5:avs_0_rmap_read_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_byteenable                  : std_logic_vector(3 downto 0);   -- mm_interconnect_1:rmap_mem_nfee_comm_5_avalon_rmap_slave_0_byteenable -> rmap_mem_nfee_comm_5:avs_0_rmap_byteenable_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_write                       : std_logic;                      -- mm_interconnect_1:rmap_mem_nfee_comm_5_avalon_rmap_slave_0_write -> rmap_mem_nfee_comm_5:avs_0_rmap_write_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:rmap_mem_nfee_comm_5_avalon_rmap_slave_0_writedata -> rmap_mem_nfee_comm_5:avs_0_rmap_writedata_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_readdata                    : std_logic_vector(31 downto 0);  -- rmap_mem_nfee_comm_6:avs_0_rmap_readdata_o -> mm_interconnect_1:rmap_mem_nfee_comm_6_avalon_rmap_slave_0_readdata
	signal mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_waitrequest                 : std_logic;                      -- rmap_mem_nfee_comm_6:avs_0_rmap_waitrequest_o -> mm_interconnect_1:rmap_mem_nfee_comm_6_avalon_rmap_slave_0_waitrequest
	signal mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_address                     : std_logic_vector(11 downto 0);  -- mm_interconnect_1:rmap_mem_nfee_comm_6_avalon_rmap_slave_0_address -> rmap_mem_nfee_comm_6:avs_0_rmap_address_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_read                        : std_logic;                      -- mm_interconnect_1:rmap_mem_nfee_comm_6_avalon_rmap_slave_0_read -> rmap_mem_nfee_comm_6:avs_0_rmap_read_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_byteenable                  : std_logic_vector(3 downto 0);   -- mm_interconnect_1:rmap_mem_nfee_comm_6_avalon_rmap_slave_0_byteenable -> rmap_mem_nfee_comm_6:avs_0_rmap_byteenable_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_write                       : std_logic;                      -- mm_interconnect_1:rmap_mem_nfee_comm_6_avalon_rmap_slave_0_write -> rmap_mem_nfee_comm_6:avs_0_rmap_write_i
	signal mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:rmap_mem_nfee_comm_6_avalon_rmap_slave_0_writedata -> rmap_mem_nfee_comm_6:avs_0_rmap_writedata_i
	signal mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_readdata                             : std_logic_vector(31 downto 0);  -- FTDI_USB3_0:avalon_slave_config_readdata -> mm_interconnect_1:FTDI_USB3_0_avalon_slave_config_readdata
	signal mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_waitrequest                          : std_logic;                      -- FTDI_USB3_0:avalon_slave_config_waitrequest -> mm_interconnect_1:FTDI_USB3_0_avalon_slave_config_waitrequest
	signal mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_address                              : std_logic_vector(7 downto 0);   -- mm_interconnect_1:FTDI_USB3_0_avalon_slave_config_address -> FTDI_USB3_0:avalon_slave_config_address
	signal mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_read                                 : std_logic;                      -- mm_interconnect_1:FTDI_USB3_0_avalon_slave_config_read -> FTDI_USB3_0:avalon_slave_config_read
	signal mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_byteenable                           : std_logic_vector(3 downto 0);   -- mm_interconnect_1:FTDI_USB3_0_avalon_slave_config_byteenable -> FTDI_USB3_0:avalon_slave_config_byteenable
	signal mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_write                                : std_logic;                      -- mm_interconnect_1:FTDI_USB3_0_avalon_slave_config_write -> FTDI_USB3_0:avalon_slave_config_write
	signal mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_writedata                            : std_logic_vector(31 downto 0);  -- mm_interconnect_1:FTDI_USB3_0_avalon_slave_config_writedata -> FTDI_USB3_0:avalon_slave_config_writedata
	signal mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_readdata                : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_A:avalon_slave_windowing_readdata -> mm_interconnect_1:COMM_Pedreiro_v1_01_A_avalon_slave_windowing_readdata
	signal mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_waitrequest             : std_logic;                      -- COMM_Pedreiro_v1_01_A:avalon_slave_windowing_waitrequest -> mm_interconnect_1:COMM_Pedreiro_v1_01_A_avalon_slave_windowing_waitrequest
	signal mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_address                 : std_logic_vector(7 downto 0);   -- mm_interconnect_1:COMM_Pedreiro_v1_01_A_avalon_slave_windowing_address -> COMM_Pedreiro_v1_01_A:avalon_slave_windowing_address
	signal mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_read                    : std_logic;                      -- mm_interconnect_1:COMM_Pedreiro_v1_01_A_avalon_slave_windowing_read -> COMM_Pedreiro_v1_01_A:avalon_slave_windowing_read
	signal mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_byteenable              : std_logic_vector(3 downto 0);   -- mm_interconnect_1:COMM_Pedreiro_v1_01_A_avalon_slave_windowing_byteenable -> COMM_Pedreiro_v1_01_A:avalon_slave_windowing_byteenable
	signal mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_write                   : std_logic;                      -- mm_interconnect_1:COMM_Pedreiro_v1_01_A_avalon_slave_windowing_write -> COMM_Pedreiro_v1_01_A:avalon_slave_windowing_write
	signal mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:COMM_Pedreiro_v1_01_A_avalon_slave_windowing_writedata -> COMM_Pedreiro_v1_01_A:avalon_slave_windowing_writedata
	signal mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_readdata                : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_B:avalon_slave_windowing_readdata -> mm_interconnect_1:COMM_Pedreiro_v1_01_B_avalon_slave_windowing_readdata
	signal mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_waitrequest             : std_logic;                      -- COMM_Pedreiro_v1_01_B:avalon_slave_windowing_waitrequest -> mm_interconnect_1:COMM_Pedreiro_v1_01_B_avalon_slave_windowing_waitrequest
	signal mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_address                 : std_logic_vector(7 downto 0);   -- mm_interconnect_1:COMM_Pedreiro_v1_01_B_avalon_slave_windowing_address -> COMM_Pedreiro_v1_01_B:avalon_slave_windowing_address
	signal mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_read                    : std_logic;                      -- mm_interconnect_1:COMM_Pedreiro_v1_01_B_avalon_slave_windowing_read -> COMM_Pedreiro_v1_01_B:avalon_slave_windowing_read
	signal mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_byteenable              : std_logic_vector(3 downto 0);   -- mm_interconnect_1:COMM_Pedreiro_v1_01_B_avalon_slave_windowing_byteenable -> COMM_Pedreiro_v1_01_B:avalon_slave_windowing_byteenable
	signal mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_write                   : std_logic;                      -- mm_interconnect_1:COMM_Pedreiro_v1_01_B_avalon_slave_windowing_write -> COMM_Pedreiro_v1_01_B:avalon_slave_windowing_write
	signal mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:COMM_Pedreiro_v1_01_B_avalon_slave_windowing_writedata -> COMM_Pedreiro_v1_01_B:avalon_slave_windowing_writedata
	signal mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_readdata                : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_C:avalon_slave_windowing_readdata -> mm_interconnect_1:COMM_Pedreiro_v1_01_C_avalon_slave_windowing_readdata
	signal mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_waitrequest             : std_logic;                      -- COMM_Pedreiro_v1_01_C:avalon_slave_windowing_waitrequest -> mm_interconnect_1:COMM_Pedreiro_v1_01_C_avalon_slave_windowing_waitrequest
	signal mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_address                 : std_logic_vector(7 downto 0);   -- mm_interconnect_1:COMM_Pedreiro_v1_01_C_avalon_slave_windowing_address -> COMM_Pedreiro_v1_01_C:avalon_slave_windowing_address
	signal mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_read                    : std_logic;                      -- mm_interconnect_1:COMM_Pedreiro_v1_01_C_avalon_slave_windowing_read -> COMM_Pedreiro_v1_01_C:avalon_slave_windowing_read
	signal mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_byteenable              : std_logic_vector(3 downto 0);   -- mm_interconnect_1:COMM_Pedreiro_v1_01_C_avalon_slave_windowing_byteenable -> COMM_Pedreiro_v1_01_C:avalon_slave_windowing_byteenable
	signal mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_write                   : std_logic;                      -- mm_interconnect_1:COMM_Pedreiro_v1_01_C_avalon_slave_windowing_write -> COMM_Pedreiro_v1_01_C:avalon_slave_windowing_write
	signal mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:COMM_Pedreiro_v1_01_C_avalon_slave_windowing_writedata -> COMM_Pedreiro_v1_01_C:avalon_slave_windowing_writedata
	signal mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_readdata                : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_D:avalon_slave_windowing_readdata -> mm_interconnect_1:COMM_Pedreiro_v1_01_D_avalon_slave_windowing_readdata
	signal mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_waitrequest             : std_logic;                      -- COMM_Pedreiro_v1_01_D:avalon_slave_windowing_waitrequest -> mm_interconnect_1:COMM_Pedreiro_v1_01_D_avalon_slave_windowing_waitrequest
	signal mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_address                 : std_logic_vector(7 downto 0);   -- mm_interconnect_1:COMM_Pedreiro_v1_01_D_avalon_slave_windowing_address -> COMM_Pedreiro_v1_01_D:avalon_slave_windowing_address
	signal mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_read                    : std_logic;                      -- mm_interconnect_1:COMM_Pedreiro_v1_01_D_avalon_slave_windowing_read -> COMM_Pedreiro_v1_01_D:avalon_slave_windowing_read
	signal mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_byteenable              : std_logic_vector(3 downto 0);   -- mm_interconnect_1:COMM_Pedreiro_v1_01_D_avalon_slave_windowing_byteenable -> COMM_Pedreiro_v1_01_D:avalon_slave_windowing_byteenable
	signal mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_write                   : std_logic;                      -- mm_interconnect_1:COMM_Pedreiro_v1_01_D_avalon_slave_windowing_write -> COMM_Pedreiro_v1_01_D:avalon_slave_windowing_write
	signal mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:COMM_Pedreiro_v1_01_D_avalon_slave_windowing_writedata -> COMM_Pedreiro_v1_01_D:avalon_slave_windowing_writedata
	signal mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_readdata                : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_E:avalon_slave_windowing_readdata -> mm_interconnect_1:COMM_Pedreiro_v1_01_E_avalon_slave_windowing_readdata
	signal mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_waitrequest             : std_logic;                      -- COMM_Pedreiro_v1_01_E:avalon_slave_windowing_waitrequest -> mm_interconnect_1:COMM_Pedreiro_v1_01_E_avalon_slave_windowing_waitrequest
	signal mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_address                 : std_logic_vector(7 downto 0);   -- mm_interconnect_1:COMM_Pedreiro_v1_01_E_avalon_slave_windowing_address -> COMM_Pedreiro_v1_01_E:avalon_slave_windowing_address
	signal mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_read                    : std_logic;                      -- mm_interconnect_1:COMM_Pedreiro_v1_01_E_avalon_slave_windowing_read -> COMM_Pedreiro_v1_01_E:avalon_slave_windowing_read
	signal mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_byteenable              : std_logic_vector(3 downto 0);   -- mm_interconnect_1:COMM_Pedreiro_v1_01_E_avalon_slave_windowing_byteenable -> COMM_Pedreiro_v1_01_E:avalon_slave_windowing_byteenable
	signal mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_write                   : std_logic;                      -- mm_interconnect_1:COMM_Pedreiro_v1_01_E_avalon_slave_windowing_write -> COMM_Pedreiro_v1_01_E:avalon_slave_windowing_write
	signal mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:COMM_Pedreiro_v1_01_E_avalon_slave_windowing_writedata -> COMM_Pedreiro_v1_01_E:avalon_slave_windowing_writedata
	signal mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_readdata                : std_logic_vector(31 downto 0);  -- COMM_Pedreiro_v1_01_F:avalon_slave_windowing_readdata -> mm_interconnect_1:COMM_Pedreiro_v1_01_F_avalon_slave_windowing_readdata
	signal mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_waitrequest             : std_logic;                      -- COMM_Pedreiro_v1_01_F:avalon_slave_windowing_waitrequest -> mm_interconnect_1:COMM_Pedreiro_v1_01_F_avalon_slave_windowing_waitrequest
	signal mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_address                 : std_logic_vector(7 downto 0);   -- mm_interconnect_1:COMM_Pedreiro_v1_01_F_avalon_slave_windowing_address -> COMM_Pedreiro_v1_01_F:avalon_slave_windowing_address
	signal mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_read                    : std_logic;                      -- mm_interconnect_1:COMM_Pedreiro_v1_01_F_avalon_slave_windowing_read -> COMM_Pedreiro_v1_01_F:avalon_slave_windowing_read
	signal mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_byteenable              : std_logic_vector(3 downto 0);   -- mm_interconnect_1:COMM_Pedreiro_v1_01_F_avalon_slave_windowing_byteenable -> COMM_Pedreiro_v1_01_F:avalon_slave_windowing_byteenable
	signal mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_write                   : std_logic;                      -- mm_interconnect_1:COMM_Pedreiro_v1_01_F_avalon_slave_windowing_write -> COMM_Pedreiro_v1_01_F:avalon_slave_windowing_write
	signal mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:COMM_Pedreiro_v1_01_F_avalon_slave_windowing_writedata -> COMM_Pedreiro_v1_01_F:avalon_slave_windowing_writedata
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_readdata                             : std_logic_vector(63 downto 0);  -- ddr2_address_span_extender:avs_cntl_readdata -> mm_interconnect_1:ddr2_address_span_extender_cntl_readdata
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_read                                 : std_logic;                      -- mm_interconnect_1:ddr2_address_span_extender_cntl_read -> ddr2_address_span_extender:avs_cntl_read
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_byteenable                           : std_logic_vector(7 downto 0);   -- mm_interconnect_1:ddr2_address_span_extender_cntl_byteenable -> ddr2_address_span_extender:avs_cntl_byteenable
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_write                                : std_logic;                      -- mm_interconnect_1:ddr2_address_span_extender_cntl_write -> ddr2_address_span_extender:avs_cntl_write
	signal mm_interconnect_1_ddr2_address_span_extender_cntl_writedata                            : std_logic_vector(63 downto 0);  -- mm_interconnect_1:ddr2_address_span_extender_cntl_writedata -> ddr2_address_span_extender:avs_cntl_writedata
	signal mm_interconnect_1_sysid_qsys_control_slave_readdata                                    : std_logic_vector(31 downto 0);  -- sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	signal mm_interconnect_1_sysid_qsys_control_slave_address                                     : std_logic_vector(0 downto 0);   -- mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	signal mm_interconnect_1_dma_comm_1_left_csr_readdata                                         : std_logic_vector(31 downto 0);  -- dma_comm_1_left:csr_readdata -> mm_interconnect_1:dma_comm_1_left_csr_readdata
	signal mm_interconnect_1_dma_comm_1_left_csr_address                                          : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_comm_1_left_csr_address -> dma_comm_1_left:csr_address
	signal mm_interconnect_1_dma_comm_1_left_csr_read                                             : std_logic;                      -- mm_interconnect_1:dma_comm_1_left_csr_read -> dma_comm_1_left:csr_read
	signal mm_interconnect_1_dma_comm_1_left_csr_byteenable                                       : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_comm_1_left_csr_byteenable -> dma_comm_1_left:csr_byteenable
	signal mm_interconnect_1_dma_comm_1_left_csr_write                                            : std_logic;                      -- mm_interconnect_1:dma_comm_1_left_csr_write -> dma_comm_1_left:csr_write
	signal mm_interconnect_1_dma_comm_1_left_csr_writedata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_1_left_csr_writedata -> dma_comm_1_left:csr_writedata
	signal mm_interconnect_1_dma_comm_1_right_csr_readdata                                        : std_logic_vector(31 downto 0);  -- dma_comm_1_right:csr_readdata -> mm_interconnect_1:dma_comm_1_right_csr_readdata
	signal mm_interconnect_1_dma_comm_1_right_csr_address                                         : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_comm_1_right_csr_address -> dma_comm_1_right:csr_address
	signal mm_interconnect_1_dma_comm_1_right_csr_read                                            : std_logic;                      -- mm_interconnect_1:dma_comm_1_right_csr_read -> dma_comm_1_right:csr_read
	signal mm_interconnect_1_dma_comm_1_right_csr_byteenable                                      : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_comm_1_right_csr_byteenable -> dma_comm_1_right:csr_byteenable
	signal mm_interconnect_1_dma_comm_1_right_csr_write                                           : std_logic;                      -- mm_interconnect_1:dma_comm_1_right_csr_write -> dma_comm_1_right:csr_write
	signal mm_interconnect_1_dma_comm_1_right_csr_writedata                                       : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_1_right_csr_writedata -> dma_comm_1_right:csr_writedata
	signal mm_interconnect_1_dma_comm_2_left_csr_readdata                                         : std_logic_vector(31 downto 0);  -- dma_comm_2_left:csr_readdata -> mm_interconnect_1:dma_comm_2_left_csr_readdata
	signal mm_interconnect_1_dma_comm_2_left_csr_address                                          : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_comm_2_left_csr_address -> dma_comm_2_left:csr_address
	signal mm_interconnect_1_dma_comm_2_left_csr_read                                             : std_logic;                      -- mm_interconnect_1:dma_comm_2_left_csr_read -> dma_comm_2_left:csr_read
	signal mm_interconnect_1_dma_comm_2_left_csr_byteenable                                       : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_comm_2_left_csr_byteenable -> dma_comm_2_left:csr_byteenable
	signal mm_interconnect_1_dma_comm_2_left_csr_write                                            : std_logic;                      -- mm_interconnect_1:dma_comm_2_left_csr_write -> dma_comm_2_left:csr_write
	signal mm_interconnect_1_dma_comm_2_left_csr_writedata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_2_left_csr_writedata -> dma_comm_2_left:csr_writedata
	signal mm_interconnect_1_dma_comm_2_right_csr_readdata                                        : std_logic_vector(31 downto 0);  -- dma_comm_2_right:csr_readdata -> mm_interconnect_1:dma_comm_2_right_csr_readdata
	signal mm_interconnect_1_dma_comm_2_right_csr_address                                         : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_comm_2_right_csr_address -> dma_comm_2_right:csr_address
	signal mm_interconnect_1_dma_comm_2_right_csr_read                                            : std_logic;                      -- mm_interconnect_1:dma_comm_2_right_csr_read -> dma_comm_2_right:csr_read
	signal mm_interconnect_1_dma_comm_2_right_csr_byteenable                                      : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_comm_2_right_csr_byteenable -> dma_comm_2_right:csr_byteenable
	signal mm_interconnect_1_dma_comm_2_right_csr_write                                           : std_logic;                      -- mm_interconnect_1:dma_comm_2_right_csr_write -> dma_comm_2_right:csr_write
	signal mm_interconnect_1_dma_comm_2_right_csr_writedata                                       : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_2_right_csr_writedata -> dma_comm_2_right:csr_writedata
	signal mm_interconnect_1_dma_comm_3_left_csr_readdata                                         : std_logic_vector(31 downto 0);  -- dma_comm_3_left:csr_readdata -> mm_interconnect_1:dma_comm_3_left_csr_readdata
	signal mm_interconnect_1_dma_comm_3_left_csr_address                                          : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_comm_3_left_csr_address -> dma_comm_3_left:csr_address
	signal mm_interconnect_1_dma_comm_3_left_csr_read                                             : std_logic;                      -- mm_interconnect_1:dma_comm_3_left_csr_read -> dma_comm_3_left:csr_read
	signal mm_interconnect_1_dma_comm_3_left_csr_byteenable                                       : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_comm_3_left_csr_byteenable -> dma_comm_3_left:csr_byteenable
	signal mm_interconnect_1_dma_comm_3_left_csr_write                                            : std_logic;                      -- mm_interconnect_1:dma_comm_3_left_csr_write -> dma_comm_3_left:csr_write
	signal mm_interconnect_1_dma_comm_3_left_csr_writedata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_3_left_csr_writedata -> dma_comm_3_left:csr_writedata
	signal mm_interconnect_1_dma_comm_3_right_csr_readdata                                        : std_logic_vector(31 downto 0);  -- dma_comm_3_right:csr_readdata -> mm_interconnect_1:dma_comm_3_right_csr_readdata
	signal mm_interconnect_1_dma_comm_3_right_csr_address                                         : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_comm_3_right_csr_address -> dma_comm_3_right:csr_address
	signal mm_interconnect_1_dma_comm_3_right_csr_read                                            : std_logic;                      -- mm_interconnect_1:dma_comm_3_right_csr_read -> dma_comm_3_right:csr_read
	signal mm_interconnect_1_dma_comm_3_right_csr_byteenable                                      : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_comm_3_right_csr_byteenable -> dma_comm_3_right:csr_byteenable
	signal mm_interconnect_1_dma_comm_3_right_csr_write                                           : std_logic;                      -- mm_interconnect_1:dma_comm_3_right_csr_write -> dma_comm_3_right:csr_write
	signal mm_interconnect_1_dma_comm_3_right_csr_writedata                                       : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_3_right_csr_writedata -> dma_comm_3_right:csr_writedata
	signal mm_interconnect_1_dma_comm_4_left_csr_readdata                                         : std_logic_vector(31 downto 0);  -- dma_comm_4_left:csr_readdata -> mm_interconnect_1:dma_comm_4_left_csr_readdata
	signal mm_interconnect_1_dma_comm_4_left_csr_address                                          : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_comm_4_left_csr_address -> dma_comm_4_left:csr_address
	signal mm_interconnect_1_dma_comm_4_left_csr_read                                             : std_logic;                      -- mm_interconnect_1:dma_comm_4_left_csr_read -> dma_comm_4_left:csr_read
	signal mm_interconnect_1_dma_comm_4_left_csr_byteenable                                       : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_comm_4_left_csr_byteenable -> dma_comm_4_left:csr_byteenable
	signal mm_interconnect_1_dma_comm_4_left_csr_write                                            : std_logic;                      -- mm_interconnect_1:dma_comm_4_left_csr_write -> dma_comm_4_left:csr_write
	signal mm_interconnect_1_dma_comm_4_left_csr_writedata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_4_left_csr_writedata -> dma_comm_4_left:csr_writedata
	signal mm_interconnect_1_dma_comm_4_right_csr_readdata                                        : std_logic_vector(31 downto 0);  -- dma_comm_4_right:csr_readdata -> mm_interconnect_1:dma_comm_4_right_csr_readdata
	signal mm_interconnect_1_dma_comm_4_right_csr_address                                         : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_comm_4_right_csr_address -> dma_comm_4_right:csr_address
	signal mm_interconnect_1_dma_comm_4_right_csr_read                                            : std_logic;                      -- mm_interconnect_1:dma_comm_4_right_csr_read -> dma_comm_4_right:csr_read
	signal mm_interconnect_1_dma_comm_4_right_csr_byteenable                                      : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_comm_4_right_csr_byteenable -> dma_comm_4_right:csr_byteenable
	signal mm_interconnect_1_dma_comm_4_right_csr_write                                           : std_logic;                      -- mm_interconnect_1:dma_comm_4_right_csr_write -> dma_comm_4_right:csr_write
	signal mm_interconnect_1_dma_comm_4_right_csr_writedata                                       : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_4_right_csr_writedata -> dma_comm_4_right:csr_writedata
	signal mm_interconnect_1_dma_comm_5_left_csr_readdata                                         : std_logic_vector(31 downto 0);  -- dma_comm_5_left:csr_readdata -> mm_interconnect_1:dma_comm_5_left_csr_readdata
	signal mm_interconnect_1_dma_comm_5_left_csr_address                                          : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_comm_5_left_csr_address -> dma_comm_5_left:csr_address
	signal mm_interconnect_1_dma_comm_5_left_csr_read                                             : std_logic;                      -- mm_interconnect_1:dma_comm_5_left_csr_read -> dma_comm_5_left:csr_read
	signal mm_interconnect_1_dma_comm_5_left_csr_byteenable                                       : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_comm_5_left_csr_byteenable -> dma_comm_5_left:csr_byteenable
	signal mm_interconnect_1_dma_comm_5_left_csr_write                                            : std_logic;                      -- mm_interconnect_1:dma_comm_5_left_csr_write -> dma_comm_5_left:csr_write
	signal mm_interconnect_1_dma_comm_5_left_csr_writedata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_5_left_csr_writedata -> dma_comm_5_left:csr_writedata
	signal mm_interconnect_1_dma_comm_5_right_csr_readdata                                        : std_logic_vector(31 downto 0);  -- dma_comm_5_right:csr_readdata -> mm_interconnect_1:dma_comm_5_right_csr_readdata
	signal mm_interconnect_1_dma_comm_5_right_csr_address                                         : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_comm_5_right_csr_address -> dma_comm_5_right:csr_address
	signal mm_interconnect_1_dma_comm_5_right_csr_read                                            : std_logic;                      -- mm_interconnect_1:dma_comm_5_right_csr_read -> dma_comm_5_right:csr_read
	signal mm_interconnect_1_dma_comm_5_right_csr_byteenable                                      : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_comm_5_right_csr_byteenable -> dma_comm_5_right:csr_byteenable
	signal mm_interconnect_1_dma_comm_5_right_csr_write                                           : std_logic;                      -- mm_interconnect_1:dma_comm_5_right_csr_write -> dma_comm_5_right:csr_write
	signal mm_interconnect_1_dma_comm_5_right_csr_writedata                                       : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_5_right_csr_writedata -> dma_comm_5_right:csr_writedata
	signal mm_interconnect_1_dma_comm_6_left_csr_readdata                                         : std_logic_vector(31 downto 0);  -- dma_comm_6_left:csr_readdata -> mm_interconnect_1:dma_comm_6_left_csr_readdata
	signal mm_interconnect_1_dma_comm_6_left_csr_address                                          : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_comm_6_left_csr_address -> dma_comm_6_left:csr_address
	signal mm_interconnect_1_dma_comm_6_left_csr_read                                             : std_logic;                      -- mm_interconnect_1:dma_comm_6_left_csr_read -> dma_comm_6_left:csr_read
	signal mm_interconnect_1_dma_comm_6_left_csr_byteenable                                       : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_comm_6_left_csr_byteenable -> dma_comm_6_left:csr_byteenable
	signal mm_interconnect_1_dma_comm_6_left_csr_write                                            : std_logic;                      -- mm_interconnect_1:dma_comm_6_left_csr_write -> dma_comm_6_left:csr_write
	signal mm_interconnect_1_dma_comm_6_left_csr_writedata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_6_left_csr_writedata -> dma_comm_6_left:csr_writedata
	signal mm_interconnect_1_dma_comm_6_right_csr_readdata                                        : std_logic_vector(31 downto 0);  -- dma_comm_6_right:csr_readdata -> mm_interconnect_1:dma_comm_6_right_csr_readdata
	signal mm_interconnect_1_dma_comm_6_right_csr_address                                         : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_comm_6_right_csr_address -> dma_comm_6_right:csr_address
	signal mm_interconnect_1_dma_comm_6_right_csr_read                                            : std_logic;                      -- mm_interconnect_1:dma_comm_6_right_csr_read -> dma_comm_6_right:csr_read
	signal mm_interconnect_1_dma_comm_6_right_csr_byteenable                                      : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_comm_6_right_csr_byteenable -> dma_comm_6_right:csr_byteenable
	signal mm_interconnect_1_dma_comm_6_right_csr_write                                           : std_logic;                      -- mm_interconnect_1:dma_comm_6_right_csr_write -> dma_comm_6_right:csr_write
	signal mm_interconnect_1_dma_comm_6_right_csr_writedata                                       : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_6_right_csr_writedata -> dma_comm_6_right:csr_writedata
	signal mm_interconnect_1_dma_ftdi_usb3_csr_readdata                                           : std_logic_vector(31 downto 0);  -- dma_ftdi_usb3:csr_readdata -> mm_interconnect_1:dma_ftdi_usb3_csr_readdata
	signal mm_interconnect_1_dma_ftdi_usb3_csr_address                                            : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_ftdi_usb3_csr_address -> dma_ftdi_usb3:csr_address
	signal mm_interconnect_1_dma_ftdi_usb3_csr_read                                               : std_logic;                      -- mm_interconnect_1:dma_ftdi_usb3_csr_read -> dma_ftdi_usb3:csr_read
	signal mm_interconnect_1_dma_ftdi_usb3_csr_byteenable                                         : std_logic_vector(3 downto 0);   -- mm_interconnect_1:dma_ftdi_usb3_csr_byteenable -> dma_ftdi_usb3:csr_byteenable
	signal mm_interconnect_1_dma_ftdi_usb3_csr_write                                              : std_logic;                      -- mm_interconnect_1:dma_ftdi_usb3_csr_write -> dma_ftdi_usb3:csr_write
	signal mm_interconnect_1_dma_ftdi_usb3_csr_writedata                                          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_ftdi_usb3_csr_writedata -> dma_ftdi_usb3:csr_writedata
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata                                : std_logic_vector(31 downto 0);  -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest                             : std_logic;                      -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess                             : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address                                 : std_logic_vector(8 downto 0);   -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read                                    : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable                              : std_logic_vector(3 downto 0);   -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write                                   : std_logic;                      -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata                               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_1_dma_comm_1_left_descriptor_slave_waitrequest                         : std_logic;                      -- dma_comm_1_left:descriptor_slave_waitrequest -> mm_interconnect_1:dma_comm_1_left_descriptor_slave_waitrequest
	signal mm_interconnect_1_dma_comm_1_left_descriptor_slave_byteenable                          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_1_left_descriptor_slave_byteenable -> dma_comm_1_left:descriptor_slave_byteenable
	signal mm_interconnect_1_dma_comm_1_left_descriptor_slave_write                               : std_logic;                      -- mm_interconnect_1:dma_comm_1_left_descriptor_slave_write -> dma_comm_1_left:descriptor_slave_write
	signal mm_interconnect_1_dma_comm_1_left_descriptor_slave_writedata                           : std_logic_vector(255 downto 0); -- mm_interconnect_1:dma_comm_1_left_descriptor_slave_writedata -> dma_comm_1_left:descriptor_slave_writedata
	signal mm_interconnect_1_dma_comm_1_right_descriptor_slave_waitrequest                        : std_logic;                      -- dma_comm_1_right:descriptor_slave_waitrequest -> mm_interconnect_1:dma_comm_1_right_descriptor_slave_waitrequest
	signal mm_interconnect_1_dma_comm_1_right_descriptor_slave_byteenable                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_1_right_descriptor_slave_byteenable -> dma_comm_1_right:descriptor_slave_byteenable
	signal mm_interconnect_1_dma_comm_1_right_descriptor_slave_write                              : std_logic;                      -- mm_interconnect_1:dma_comm_1_right_descriptor_slave_write -> dma_comm_1_right:descriptor_slave_write
	signal mm_interconnect_1_dma_comm_1_right_descriptor_slave_writedata                          : std_logic_vector(255 downto 0); -- mm_interconnect_1:dma_comm_1_right_descriptor_slave_writedata -> dma_comm_1_right:descriptor_slave_writedata
	signal mm_interconnect_1_dma_comm_2_left_descriptor_slave_waitrequest                         : std_logic;                      -- dma_comm_2_left:descriptor_slave_waitrequest -> mm_interconnect_1:dma_comm_2_left_descriptor_slave_waitrequest
	signal mm_interconnect_1_dma_comm_2_left_descriptor_slave_byteenable                          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_2_left_descriptor_slave_byteenable -> dma_comm_2_left:descriptor_slave_byteenable
	signal mm_interconnect_1_dma_comm_2_left_descriptor_slave_write                               : std_logic;                      -- mm_interconnect_1:dma_comm_2_left_descriptor_slave_write -> dma_comm_2_left:descriptor_slave_write
	signal mm_interconnect_1_dma_comm_2_left_descriptor_slave_writedata                           : std_logic_vector(255 downto 0); -- mm_interconnect_1:dma_comm_2_left_descriptor_slave_writedata -> dma_comm_2_left:descriptor_slave_writedata
	signal mm_interconnect_1_dma_comm_2_right_descriptor_slave_waitrequest                        : std_logic;                      -- dma_comm_2_right:descriptor_slave_waitrequest -> mm_interconnect_1:dma_comm_2_right_descriptor_slave_waitrequest
	signal mm_interconnect_1_dma_comm_2_right_descriptor_slave_byteenable                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_2_right_descriptor_slave_byteenable -> dma_comm_2_right:descriptor_slave_byteenable
	signal mm_interconnect_1_dma_comm_2_right_descriptor_slave_write                              : std_logic;                      -- mm_interconnect_1:dma_comm_2_right_descriptor_slave_write -> dma_comm_2_right:descriptor_slave_write
	signal mm_interconnect_1_dma_comm_2_right_descriptor_slave_writedata                          : std_logic_vector(255 downto 0); -- mm_interconnect_1:dma_comm_2_right_descriptor_slave_writedata -> dma_comm_2_right:descriptor_slave_writedata
	signal mm_interconnect_1_dma_comm_3_left_descriptor_slave_waitrequest                         : std_logic;                      -- dma_comm_3_left:descriptor_slave_waitrequest -> mm_interconnect_1:dma_comm_3_left_descriptor_slave_waitrequest
	signal mm_interconnect_1_dma_comm_3_left_descriptor_slave_byteenable                          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_3_left_descriptor_slave_byteenable -> dma_comm_3_left:descriptor_slave_byteenable
	signal mm_interconnect_1_dma_comm_3_left_descriptor_slave_write                               : std_logic;                      -- mm_interconnect_1:dma_comm_3_left_descriptor_slave_write -> dma_comm_3_left:descriptor_slave_write
	signal mm_interconnect_1_dma_comm_3_left_descriptor_slave_writedata                           : std_logic_vector(255 downto 0); -- mm_interconnect_1:dma_comm_3_left_descriptor_slave_writedata -> dma_comm_3_left:descriptor_slave_writedata
	signal mm_interconnect_1_dma_comm_3_right_descriptor_slave_waitrequest                        : std_logic;                      -- dma_comm_3_right:descriptor_slave_waitrequest -> mm_interconnect_1:dma_comm_3_right_descriptor_slave_waitrequest
	signal mm_interconnect_1_dma_comm_3_right_descriptor_slave_byteenable                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_3_right_descriptor_slave_byteenable -> dma_comm_3_right:descriptor_slave_byteenable
	signal mm_interconnect_1_dma_comm_3_right_descriptor_slave_write                              : std_logic;                      -- mm_interconnect_1:dma_comm_3_right_descriptor_slave_write -> dma_comm_3_right:descriptor_slave_write
	signal mm_interconnect_1_dma_comm_3_right_descriptor_slave_writedata                          : std_logic_vector(255 downto 0); -- mm_interconnect_1:dma_comm_3_right_descriptor_slave_writedata -> dma_comm_3_right:descriptor_slave_writedata
	signal mm_interconnect_1_dma_comm_4_left_descriptor_slave_waitrequest                         : std_logic;                      -- dma_comm_4_left:descriptor_slave_waitrequest -> mm_interconnect_1:dma_comm_4_left_descriptor_slave_waitrequest
	signal mm_interconnect_1_dma_comm_4_left_descriptor_slave_byteenable                          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_4_left_descriptor_slave_byteenable -> dma_comm_4_left:descriptor_slave_byteenable
	signal mm_interconnect_1_dma_comm_4_left_descriptor_slave_write                               : std_logic;                      -- mm_interconnect_1:dma_comm_4_left_descriptor_slave_write -> dma_comm_4_left:descriptor_slave_write
	signal mm_interconnect_1_dma_comm_4_left_descriptor_slave_writedata                           : std_logic_vector(255 downto 0); -- mm_interconnect_1:dma_comm_4_left_descriptor_slave_writedata -> dma_comm_4_left:descriptor_slave_writedata
	signal mm_interconnect_1_dma_comm_4_right_descriptor_slave_waitrequest                        : std_logic;                      -- dma_comm_4_right:descriptor_slave_waitrequest -> mm_interconnect_1:dma_comm_4_right_descriptor_slave_waitrequest
	signal mm_interconnect_1_dma_comm_4_right_descriptor_slave_byteenable                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_4_right_descriptor_slave_byteenable -> dma_comm_4_right:descriptor_slave_byteenable
	signal mm_interconnect_1_dma_comm_4_right_descriptor_slave_write                              : std_logic;                      -- mm_interconnect_1:dma_comm_4_right_descriptor_slave_write -> dma_comm_4_right:descriptor_slave_write
	signal mm_interconnect_1_dma_comm_4_right_descriptor_slave_writedata                          : std_logic_vector(255 downto 0); -- mm_interconnect_1:dma_comm_4_right_descriptor_slave_writedata -> dma_comm_4_right:descriptor_slave_writedata
	signal mm_interconnect_1_dma_comm_5_left_descriptor_slave_waitrequest                         : std_logic;                      -- dma_comm_5_left:descriptor_slave_waitrequest -> mm_interconnect_1:dma_comm_5_left_descriptor_slave_waitrequest
	signal mm_interconnect_1_dma_comm_5_left_descriptor_slave_byteenable                          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_5_left_descriptor_slave_byteenable -> dma_comm_5_left:descriptor_slave_byteenable
	signal mm_interconnect_1_dma_comm_5_left_descriptor_slave_write                               : std_logic;                      -- mm_interconnect_1:dma_comm_5_left_descriptor_slave_write -> dma_comm_5_left:descriptor_slave_write
	signal mm_interconnect_1_dma_comm_5_left_descriptor_slave_writedata                           : std_logic_vector(255 downto 0); -- mm_interconnect_1:dma_comm_5_left_descriptor_slave_writedata -> dma_comm_5_left:descriptor_slave_writedata
	signal mm_interconnect_1_dma_comm_5_right_descriptor_slave_waitrequest                        : std_logic;                      -- dma_comm_5_right:descriptor_slave_waitrequest -> mm_interconnect_1:dma_comm_5_right_descriptor_slave_waitrequest
	signal mm_interconnect_1_dma_comm_5_right_descriptor_slave_byteenable                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_5_right_descriptor_slave_byteenable -> dma_comm_5_right:descriptor_slave_byteenable
	signal mm_interconnect_1_dma_comm_5_right_descriptor_slave_write                              : std_logic;                      -- mm_interconnect_1:dma_comm_5_right_descriptor_slave_write -> dma_comm_5_right:descriptor_slave_write
	signal mm_interconnect_1_dma_comm_5_right_descriptor_slave_writedata                          : std_logic_vector(255 downto 0); -- mm_interconnect_1:dma_comm_5_right_descriptor_slave_writedata -> dma_comm_5_right:descriptor_slave_writedata
	signal mm_interconnect_1_dma_comm_6_left_descriptor_slave_waitrequest                         : std_logic;                      -- dma_comm_6_left:descriptor_slave_waitrequest -> mm_interconnect_1:dma_comm_6_left_descriptor_slave_waitrequest
	signal mm_interconnect_1_dma_comm_6_left_descriptor_slave_byteenable                          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_6_left_descriptor_slave_byteenable -> dma_comm_6_left:descriptor_slave_byteenable
	signal mm_interconnect_1_dma_comm_6_left_descriptor_slave_write                               : std_logic;                      -- mm_interconnect_1:dma_comm_6_left_descriptor_slave_write -> dma_comm_6_left:descriptor_slave_write
	signal mm_interconnect_1_dma_comm_6_left_descriptor_slave_writedata                           : std_logic_vector(255 downto 0); -- mm_interconnect_1:dma_comm_6_left_descriptor_slave_writedata -> dma_comm_6_left:descriptor_slave_writedata
	signal mm_interconnect_1_dma_comm_6_right_descriptor_slave_waitrequest                        : std_logic;                      -- dma_comm_6_right:descriptor_slave_waitrequest -> mm_interconnect_1:dma_comm_6_right_descriptor_slave_waitrequest
	signal mm_interconnect_1_dma_comm_6_right_descriptor_slave_byteenable                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_comm_6_right_descriptor_slave_byteenable -> dma_comm_6_right:descriptor_slave_byteenable
	signal mm_interconnect_1_dma_comm_6_right_descriptor_slave_write                              : std_logic;                      -- mm_interconnect_1:dma_comm_6_right_descriptor_slave_write -> dma_comm_6_right:descriptor_slave_write
	signal mm_interconnect_1_dma_comm_6_right_descriptor_slave_writedata                          : std_logic_vector(255 downto 0); -- mm_interconnect_1:dma_comm_6_right_descriptor_slave_writedata -> dma_comm_6_right:descriptor_slave_writedata
	signal mm_interconnect_1_dma_ftdi_usb3_descriptor_slave_waitrequest                           : std_logic;                      -- dma_ftdi_usb3:descriptor_slave_waitrequest -> mm_interconnect_1:dma_ftdi_usb3_descriptor_slave_waitrequest
	signal mm_interconnect_1_dma_ftdi_usb3_descriptor_slave_byteenable                            : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_ftdi_usb3_descriptor_slave_byteenable -> dma_ftdi_usb3:descriptor_slave_byteenable
	signal mm_interconnect_1_dma_ftdi_usb3_descriptor_slave_write                                 : std_logic;                      -- mm_interconnect_1:dma_ftdi_usb3_descriptor_slave_write -> dma_ftdi_usb3:descriptor_slave_write
	signal mm_interconnect_1_dma_ftdi_usb3_descriptor_slave_writedata                             : std_logic_vector(255 downto 0); -- mm_interconnect_1:dma_ftdi_usb3_descriptor_slave_writedata -> dma_ftdi_usb3:descriptor_slave_writedata
	signal mm_interconnect_1_clock_bridge_afi_50_s0_readdata                                      : std_logic_vector(31 downto 0);  -- clock_bridge_afi_50:s0_readdata -> mm_interconnect_1:clock_bridge_afi_50_s0_readdata
	signal mm_interconnect_1_clock_bridge_afi_50_s0_waitrequest                                   : std_logic;                      -- clock_bridge_afi_50:s0_waitrequest -> mm_interconnect_1:clock_bridge_afi_50_s0_waitrequest
	signal mm_interconnect_1_clock_bridge_afi_50_s0_debugaccess                                   : std_logic;                      -- mm_interconnect_1:clock_bridge_afi_50_s0_debugaccess -> clock_bridge_afi_50:s0_debugaccess
	signal mm_interconnect_1_clock_bridge_afi_50_s0_address                                       : std_logic_vector(11 downto 0);  -- mm_interconnect_1:clock_bridge_afi_50_s0_address -> clock_bridge_afi_50:s0_address
	signal mm_interconnect_1_clock_bridge_afi_50_s0_read                                          : std_logic;                      -- mm_interconnect_1:clock_bridge_afi_50_s0_read -> clock_bridge_afi_50:s0_read
	signal mm_interconnect_1_clock_bridge_afi_50_s0_byteenable                                    : std_logic_vector(3 downto 0);   -- mm_interconnect_1:clock_bridge_afi_50_s0_byteenable -> clock_bridge_afi_50:s0_byteenable
	signal mm_interconnect_1_clock_bridge_afi_50_s0_readdatavalid                                 : std_logic;                      -- clock_bridge_afi_50:s0_readdatavalid -> mm_interconnect_1:clock_bridge_afi_50_s0_readdatavalid
	signal mm_interconnect_1_clock_bridge_afi_50_s0_write                                         : std_logic;                      -- mm_interconnect_1:clock_bridge_afi_50_s0_write -> clock_bridge_afi_50:s0_write
	signal mm_interconnect_1_clock_bridge_afi_50_s0_writedata                                     : std_logic_vector(31 downto 0);  -- mm_interconnect_1:clock_bridge_afi_50_s0_writedata -> clock_bridge_afi_50:s0_writedata
	signal mm_interconnect_1_clock_bridge_afi_50_s0_burstcount                                    : std_logic_vector(0 downto 0);   -- mm_interconnect_1:clock_bridge_afi_50_s0_burstcount -> clock_bridge_afi_50:s0_burstcount
	signal mm_interconnect_1_onchip_memory_s1_chipselect                                          : std_logic;                      -- mm_interconnect_1:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	signal mm_interconnect_1_onchip_memory_s1_readdata                                            : std_logic_vector(31 downto 0);  -- onchip_memory:readdata -> mm_interconnect_1:onchip_memory_s1_readdata
	signal mm_interconnect_1_onchip_memory_s1_address                                             : std_logic_vector(17 downto 0);  -- mm_interconnect_1:onchip_memory_s1_address -> onchip_memory:address
	signal mm_interconnect_1_onchip_memory_s1_byteenable                                          : std_logic_vector(3 downto 0);   -- mm_interconnect_1:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	signal mm_interconnect_1_onchip_memory_s1_write                                               : std_logic;                      -- mm_interconnect_1:onchip_memory_s1_write -> onchip_memory:write
	signal mm_interconnect_1_onchip_memory_s1_writedata                                           : std_logic_vector(31 downto 0);  -- mm_interconnect_1:onchip_memory_s1_writedata -> onchip_memory:writedata
	signal mm_interconnect_1_onchip_memory_s1_clken                                               : std_logic;                      -- mm_interconnect_1:onchip_memory_s1_clken -> onchip_memory:clken
	signal mm_interconnect_1_ext_flash_uas_readdata                                               : std_logic_vector(15 downto 0);  -- ext_flash:uas_readdata -> mm_interconnect_1:ext_flash_uas_readdata
	signal mm_interconnect_1_ext_flash_uas_waitrequest                                            : std_logic;                      -- ext_flash:uas_waitrequest -> mm_interconnect_1:ext_flash_uas_waitrequest
	signal mm_interconnect_1_ext_flash_uas_debugaccess                                            : std_logic;                      -- mm_interconnect_1:ext_flash_uas_debugaccess -> ext_flash:uas_debugaccess
	signal mm_interconnect_1_ext_flash_uas_address                                                : std_logic_vector(25 downto 0);  -- mm_interconnect_1:ext_flash_uas_address -> ext_flash:uas_address
	signal mm_interconnect_1_ext_flash_uas_read                                                   : std_logic;                      -- mm_interconnect_1:ext_flash_uas_read -> ext_flash:uas_read
	signal mm_interconnect_1_ext_flash_uas_byteenable                                             : std_logic_vector(1 downto 0);   -- mm_interconnect_1:ext_flash_uas_byteenable -> ext_flash:uas_byteenable
	signal mm_interconnect_1_ext_flash_uas_readdatavalid                                          : std_logic;                      -- ext_flash:uas_readdatavalid -> mm_interconnect_1:ext_flash_uas_readdatavalid
	signal mm_interconnect_1_ext_flash_uas_lock                                                   : std_logic;                      -- mm_interconnect_1:ext_flash_uas_lock -> ext_flash:uas_lock
	signal mm_interconnect_1_ext_flash_uas_write                                                  : std_logic;                      -- mm_interconnect_1:ext_flash_uas_write -> ext_flash:uas_write
	signal mm_interconnect_1_ext_flash_uas_writedata                                              : std_logic_vector(15 downto 0);  -- mm_interconnect_1:ext_flash_uas_writedata -> ext_flash:uas_writedata
	signal mm_interconnect_1_ext_flash_uas_burstcount                                             : std_logic_vector(1 downto 0);   -- mm_interconnect_1:ext_flash_uas_burstcount -> ext_flash:uas_burstcount
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdata                   : std_logic_vector(31 downto 0);  -- ddr2_address_span_extender:avs_s0_readdata -> mm_interconnect_1:ddr2_address_span_extender_windowed_slave_readdata
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_waitrequest                : std_logic;                      -- ddr2_address_span_extender:avs_s0_waitrequest -> mm_interconnect_1:ddr2_address_span_extender_windowed_slave_waitrequest
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_address                    : std_logic_vector(28 downto 0);  -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_address -> ddr2_address_span_extender:avs_s0_address
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_read                       : std_logic;                      -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_read -> ddr2_address_span_extender:avs_s0_read
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_byteenable                 : std_logic_vector(3 downto 0);   -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_byteenable -> ddr2_address_span_extender:avs_s0_byteenable
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdatavalid              : std_logic;                      -- ddr2_address_span_extender:avs_s0_readdatavalid -> mm_interconnect_1:ddr2_address_span_extender_windowed_slave_readdatavalid
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_write                      : std_logic;                      -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_write -> ddr2_address_span_extender:avs_s0_write
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_writedata                  : std_logic_vector(31 downto 0);  -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_writedata -> ddr2_address_span_extender:avs_s0_writedata
	signal mm_interconnect_1_ddr2_address_span_extender_windowed_slave_burstcount                 : std_logic_vector(7 downto 0);   -- mm_interconnect_1:ddr2_address_span_extender_windowed_slave_burstcount -> ddr2_address_span_extender:avs_s0_burstcount
	signal clock_bridge_afi_50_m0_waitrequest                                                     : std_logic;                      -- mm_interconnect_2:clock_bridge_afi_50_m0_waitrequest -> clock_bridge_afi_50:m0_waitrequest
	signal clock_bridge_afi_50_m0_readdata                                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_2:clock_bridge_afi_50_m0_readdata -> clock_bridge_afi_50:m0_readdata
	signal clock_bridge_afi_50_m0_debugaccess                                                     : std_logic;                      -- clock_bridge_afi_50:m0_debugaccess -> mm_interconnect_2:clock_bridge_afi_50_m0_debugaccess
	signal clock_bridge_afi_50_m0_address                                                         : std_logic_vector(11 downto 0);  -- clock_bridge_afi_50:m0_address -> mm_interconnect_2:clock_bridge_afi_50_m0_address
	signal clock_bridge_afi_50_m0_read                                                            : std_logic;                      -- clock_bridge_afi_50:m0_read -> mm_interconnect_2:clock_bridge_afi_50_m0_read
	signal clock_bridge_afi_50_m0_byteenable                                                      : std_logic_vector(3 downto 0);   -- clock_bridge_afi_50:m0_byteenable -> mm_interconnect_2:clock_bridge_afi_50_m0_byteenable
	signal clock_bridge_afi_50_m0_readdatavalid                                                   : std_logic;                      -- mm_interconnect_2:clock_bridge_afi_50_m0_readdatavalid -> clock_bridge_afi_50:m0_readdatavalid
	signal clock_bridge_afi_50_m0_writedata                                                       : std_logic_vector(31 downto 0);  -- clock_bridge_afi_50:m0_writedata -> mm_interconnect_2:clock_bridge_afi_50_m0_writedata
	signal clock_bridge_afi_50_m0_write                                                           : std_logic;                      -- clock_bridge_afi_50:m0_write -> mm_interconnect_2:clock_bridge_afi_50_m0_write
	signal clock_bridge_afi_50_m0_burstcount                                                      : std_logic_vector(0 downto 0);   -- clock_bridge_afi_50:m0_burstcount -> mm_interconnect_2:clock_bridge_afi_50_m0_burstcount
	signal mm_interconnect_2_seven_segment_controller_0_ssdp_avalon_slave_address                 : std_logic_vector(0 downto 0);   -- mm_interconnect_2:SEVEN_SEGMENT_CONTROLLER_0_SSDP_avalon_slave_address -> SEVEN_SEGMENT_CONTROLLER_0:AVALON_SLAVE_ADDRESS
	signal mm_interconnect_2_seven_segment_controller_0_ssdp_avalon_slave_write                   : std_logic;                      -- mm_interconnect_2:SEVEN_SEGMENT_CONTROLLER_0_SSDP_avalon_slave_write -> SEVEN_SEGMENT_CONTROLLER_0:AVALON_SLAVE_WRITE
	signal mm_interconnect_2_seven_segment_controller_0_ssdp_avalon_slave_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_2:SEVEN_SEGMENT_CONTROLLER_0_SSDP_avalon_slave_writedata -> SEVEN_SEGMENT_CONTROLLER_0:AVALON_SLAVE_WRITEDATA
	signal mm_interconnect_2_sync_avalon_mm_slave_readdata                                        : std_logic_vector(31 downto 0);  -- sync:avalon_slave_readdata_o -> mm_interconnect_2:sync_avalon_mm_slave_readdata
	signal mm_interconnect_2_sync_avalon_mm_slave_waitrequest                                     : std_logic;                      -- sync:avalon_slave_waitrequest_o -> mm_interconnect_2:sync_avalon_mm_slave_waitrequest
	signal mm_interconnect_2_sync_avalon_mm_slave_address                                         : std_logic_vector(7 downto 0);   -- mm_interconnect_2:sync_avalon_mm_slave_address -> sync:avalon_slave_address_i
	signal mm_interconnect_2_sync_avalon_mm_slave_read                                            : std_logic;                      -- mm_interconnect_2:sync_avalon_mm_slave_read -> sync:avalon_slave_read_i
	signal mm_interconnect_2_sync_avalon_mm_slave_byteenable                                      : std_logic_vector(3 downto 0);   -- mm_interconnect_2:sync_avalon_mm_slave_byteenable -> sync:avalon_slave_byteenable_i
	signal mm_interconnect_2_sync_avalon_mm_slave_write                                           : std_logic;                      -- mm_interconnect_2:sync_avalon_mm_slave_write -> sync:avalon_slave_write_i
	signal mm_interconnect_2_sync_avalon_mm_slave_writedata                                       : std_logic_vector(31 downto 0);  -- mm_interconnect_2:sync_avalon_mm_slave_writedata -> sync:avalon_slave_writedata_i
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_readdata                  : std_logic_vector(31 downto 0);  -- rst_controller:avalon_slave_rst_controller_readdata -> mm_interconnect_2:rst_controller_avalon_rst_controller_slave_readdata
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_waitrequest               : std_logic;                      -- rst_controller:avalon_slave_rst_controller_waitrequest -> mm_interconnect_2:rst_controller_avalon_rst_controller_slave_waitrequest
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_address                   : std_logic_vector(3 downto 0);   -- mm_interconnect_2:rst_controller_avalon_rst_controller_slave_address -> rst_controller:avalon_slave_rst_controller_address
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_read                      : std_logic;                      -- mm_interconnect_2:rst_controller_avalon_rst_controller_slave_read -> rst_controller:avalon_slave_rst_controller_read
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_write                     : std_logic;                      -- mm_interconnect_2:rst_controller_avalon_rst_controller_slave_write -> rst_controller:avalon_slave_rst_controller_write
	signal mm_interconnect_2_rst_controller_avalon_rst_controller_slave_writedata                 : std_logic_vector(31 downto 0);  -- mm_interconnect_2:rst_controller_avalon_rst_controller_slave_writedata -> rst_controller:avalon_slave_rst_controller_writedata
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect  : std_logic;                      -- mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_chip_select
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata    : std_logic_vector(31 downto 0);  -- Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_readdata -> mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest : std_logic;                      -- Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_waitrequest -> mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address     : std_logic_vector(7 downto 0);   -- mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_address
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read        : std_logic;                      -- mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_read
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable  : std_logic_vector(3 downto 0);   -- mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_byteenable
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write       : std_logic;                      -- mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_write
	signal mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata   : std_logic_vector(31 downto 0);  -- mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_writedata
	signal mm_interconnect_2_m1_ddr2_i2c_sda_s1_chipselect                                        : std_logic;                      -- mm_interconnect_2:m1_ddr2_i2c_sda_s1_chipselect -> m1_ddr2_i2c_sda:chipselect
	signal mm_interconnect_2_m1_ddr2_i2c_sda_s1_readdata                                          : std_logic_vector(31 downto 0);  -- m1_ddr2_i2c_sda:readdata -> mm_interconnect_2:m1_ddr2_i2c_sda_s1_readdata
	signal mm_interconnect_2_m1_ddr2_i2c_sda_s1_address                                           : std_logic_vector(1 downto 0);   -- mm_interconnect_2:m1_ddr2_i2c_sda_s1_address -> m1_ddr2_i2c_sda:address
	signal mm_interconnect_2_m1_ddr2_i2c_sda_s1_write                                             : std_logic;                      -- mm_interconnect_2:m1_ddr2_i2c_sda_s1_write -> mm_interconnect_2_m1_ddr2_i2c_sda_s1_write:in
	signal mm_interconnect_2_m1_ddr2_i2c_sda_s1_writedata                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_2:m1_ddr2_i2c_sda_s1_writedata -> m1_ddr2_i2c_sda:writedata
	signal mm_interconnect_2_m1_ddr2_i2c_scl_s1_chipselect                                        : std_logic;                      -- mm_interconnect_2:m1_ddr2_i2c_scl_s1_chipselect -> m1_ddr2_i2c_scl:chipselect
	signal mm_interconnect_2_m1_ddr2_i2c_scl_s1_readdata                                          : std_logic_vector(31 downto 0);  -- m1_ddr2_i2c_scl:readdata -> mm_interconnect_2:m1_ddr2_i2c_scl_s1_readdata
	signal mm_interconnect_2_m1_ddr2_i2c_scl_s1_address                                           : std_logic_vector(1 downto 0);   -- mm_interconnect_2:m1_ddr2_i2c_scl_s1_address -> m1_ddr2_i2c_scl:address
	signal mm_interconnect_2_m1_ddr2_i2c_scl_s1_write                                             : std_logic;                      -- mm_interconnect_2:m1_ddr2_i2c_scl_s1_write -> mm_interconnect_2_m1_ddr2_i2c_scl_s1_write:in
	signal mm_interconnect_2_m1_ddr2_i2c_scl_s1_writedata                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_2:m1_ddr2_i2c_scl_s1_writedata -> m1_ddr2_i2c_scl:writedata
	signal mm_interconnect_2_pio_button_s1_readdata                                               : std_logic_vector(31 downto 0);  -- pio_BUTTON:readdata -> mm_interconnect_2:pio_BUTTON_s1_readdata
	signal mm_interconnect_2_pio_button_s1_address                                                : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_BUTTON_s1_address -> pio_BUTTON:address
	signal mm_interconnect_2_pio_led_s1_chipselect                                                : std_logic;                      -- mm_interconnect_2:pio_LED_s1_chipselect -> pio_LED:chipselect
	signal mm_interconnect_2_pio_led_s1_readdata                                                  : std_logic_vector(31 downto 0);  -- pio_LED:readdata -> mm_interconnect_2:pio_LED_s1_readdata
	signal mm_interconnect_2_pio_led_s1_address                                                   : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_LED_s1_address -> pio_LED:address
	signal mm_interconnect_2_pio_led_s1_write                                                     : std_logic;                      -- mm_interconnect_2:pio_LED_s1_write -> mm_interconnect_2_pio_led_s1_write:in
	signal mm_interconnect_2_pio_led_s1_writedata                                                 : std_logic_vector(31 downto 0);  -- mm_interconnect_2:pio_LED_s1_writedata -> pio_LED:writedata
	signal mm_interconnect_2_timer_1ms_s1_chipselect                                              : std_logic;                      -- mm_interconnect_2:timer_1ms_s1_chipselect -> timer_1ms:chipselect
	signal mm_interconnect_2_timer_1ms_s1_readdata                                                : std_logic_vector(15 downto 0);  -- timer_1ms:readdata -> mm_interconnect_2:timer_1ms_s1_readdata
	signal mm_interconnect_2_timer_1ms_s1_address                                                 : std_logic_vector(2 downto 0);   -- mm_interconnect_2:timer_1ms_s1_address -> timer_1ms:address
	signal mm_interconnect_2_timer_1ms_s1_write                                                   : std_logic;                      -- mm_interconnect_2:timer_1ms_s1_write -> mm_interconnect_2_timer_1ms_s1_write:in
	signal mm_interconnect_2_timer_1ms_s1_writedata                                               : std_logic_vector(15 downto 0);  -- mm_interconnect_2:timer_1ms_s1_writedata -> timer_1ms:writedata
	signal mm_interconnect_2_pio_dip_s1_readdata                                                  : std_logic_vector(31 downto 0);  -- pio_DIP:readdata -> mm_interconnect_2:pio_DIP_s1_readdata
	signal mm_interconnect_2_pio_dip_s1_address                                                   : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_DIP_s1_address -> pio_DIP:address
	signal mm_interconnect_2_timer_1us_s1_chipselect                                              : std_logic;                      -- mm_interconnect_2:timer_1us_s1_chipselect -> timer_1us:chipselect
	signal mm_interconnect_2_timer_1us_s1_readdata                                                : std_logic_vector(15 downto 0);  -- timer_1us:readdata -> mm_interconnect_2:timer_1us_s1_readdata
	signal mm_interconnect_2_timer_1us_s1_address                                                 : std_logic_vector(2 downto 0);   -- mm_interconnect_2:timer_1us_s1_address -> timer_1us:address
	signal mm_interconnect_2_timer_1us_s1_write                                                   : std_logic;                      -- mm_interconnect_2:timer_1us_s1_write -> mm_interconnect_2_timer_1us_s1_write:in
	signal mm_interconnect_2_timer_1us_s1_writedata                                               : std_logic_vector(15 downto 0);  -- mm_interconnect_2:timer_1us_s1_writedata -> timer_1us:writedata
	signal mm_interconnect_2_pio_ext_s1_readdata                                                  : std_logic_vector(31 downto 0);  -- pio_EXT:readdata -> mm_interconnect_2:pio_EXT_s1_readdata
	signal mm_interconnect_2_pio_ext_s1_address                                                   : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_EXT_s1_address -> pio_EXT:address
	signal mm_interconnect_2_sd_card_wp_n_s1_readdata                                             : std_logic_vector(31 downto 0);  -- sd_card_wp_n:readdata -> mm_interconnect_2:sd_card_wp_n_s1_readdata
	signal mm_interconnect_2_sd_card_wp_n_s1_address                                              : std_logic_vector(1 downto 0);   -- mm_interconnect_2:sd_card_wp_n_s1_address -> sd_card_wp_n:address
	signal mm_interconnect_2_temp_scl_s1_chipselect                                               : std_logic;                      -- mm_interconnect_2:temp_scl_s1_chipselect -> temp_scl:chipselect
	signal mm_interconnect_2_temp_scl_s1_readdata                                                 : std_logic_vector(31 downto 0);  -- temp_scl:readdata -> mm_interconnect_2:temp_scl_s1_readdata
	signal mm_interconnect_2_temp_scl_s1_address                                                  : std_logic_vector(1 downto 0);   -- mm_interconnect_2:temp_scl_s1_address -> temp_scl:address
	signal mm_interconnect_2_temp_scl_s1_write                                                    : std_logic;                      -- mm_interconnect_2:temp_scl_s1_write -> mm_interconnect_2_temp_scl_s1_write:in
	signal mm_interconnect_2_temp_scl_s1_writedata                                                : std_logic_vector(31 downto 0);  -- mm_interconnect_2:temp_scl_s1_writedata -> temp_scl:writedata
	signal mm_interconnect_2_temp_sda_s1_chipselect                                               : std_logic;                      -- mm_interconnect_2:temp_sda_s1_chipselect -> temp_sda:chipselect
	signal mm_interconnect_2_temp_sda_s1_readdata                                                 : std_logic_vector(31 downto 0);  -- temp_sda:readdata -> mm_interconnect_2:temp_sda_s1_readdata
	signal mm_interconnect_2_temp_sda_s1_address                                                  : std_logic_vector(1 downto 0);   -- mm_interconnect_2:temp_sda_s1_address -> temp_sda:address
	signal mm_interconnect_2_temp_sda_s1_write                                                    : std_logic;                      -- mm_interconnect_2:temp_sda_s1_write -> mm_interconnect_2_temp_sda_s1_write:in
	signal mm_interconnect_2_temp_sda_s1_writedata                                                : std_logic_vector(31 downto 0);  -- mm_interconnect_2:temp_sda_s1_writedata -> temp_sda:writedata
	signal mm_interconnect_2_m2_ddr2_i2c_sda_s1_chipselect                                        : std_logic;                      -- mm_interconnect_2:m2_ddr2_i2c_sda_s1_chipselect -> m2_ddr2_i2c_sda:chipselect
	signal mm_interconnect_2_m2_ddr2_i2c_sda_s1_readdata                                          : std_logic_vector(31 downto 0);  -- m2_ddr2_i2c_sda:readdata -> mm_interconnect_2:m2_ddr2_i2c_sda_s1_readdata
	signal mm_interconnect_2_m2_ddr2_i2c_sda_s1_address                                           : std_logic_vector(1 downto 0);   -- mm_interconnect_2:m2_ddr2_i2c_sda_s1_address -> m2_ddr2_i2c_sda:address
	signal mm_interconnect_2_m2_ddr2_i2c_sda_s1_write                                             : std_logic;                      -- mm_interconnect_2:m2_ddr2_i2c_sda_s1_write -> mm_interconnect_2_m2_ddr2_i2c_sda_s1_write:in
	signal mm_interconnect_2_m2_ddr2_i2c_sda_s1_writedata                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_2:m2_ddr2_i2c_sda_s1_writedata -> m2_ddr2_i2c_sda:writedata
	signal mm_interconnect_2_m2_ddr2_i2c_scl_s1_chipselect                                        : std_logic;                      -- mm_interconnect_2:m2_ddr2_i2c_scl_s1_chipselect -> m2_ddr2_i2c_scl:chipselect
	signal mm_interconnect_2_m2_ddr2_i2c_scl_s1_readdata                                          : std_logic_vector(31 downto 0);  -- m2_ddr2_i2c_scl:readdata -> mm_interconnect_2:m2_ddr2_i2c_scl_s1_readdata
	signal mm_interconnect_2_m2_ddr2_i2c_scl_s1_address                                           : std_logic_vector(1 downto 0);   -- mm_interconnect_2:m2_ddr2_i2c_scl_s1_address -> m2_ddr2_i2c_scl:address
	signal mm_interconnect_2_m2_ddr2_i2c_scl_s1_write                                             : std_logic;                      -- mm_interconnect_2:m2_ddr2_i2c_scl_s1_write -> mm_interconnect_2_m2_ddr2_i2c_scl_s1_write:in
	signal mm_interconnect_2_m2_ddr2_i2c_scl_s1_writedata                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_2:m2_ddr2_i2c_scl_s1_writedata -> m2_ddr2_i2c_scl:writedata
	signal mm_interconnect_2_csense_sdo_s1_readdata                                               : std_logic_vector(31 downto 0);  -- csense_sdo:readdata -> mm_interconnect_2:csense_sdo_s1_readdata
	signal mm_interconnect_2_csense_sdo_s1_address                                                : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_sdo_s1_address -> csense_sdo:address
	signal mm_interconnect_2_csense_sdi_s1_chipselect                                             : std_logic;                      -- mm_interconnect_2:csense_sdi_s1_chipselect -> csense_sdi:chipselect
	signal mm_interconnect_2_csense_sdi_s1_readdata                                               : std_logic_vector(31 downto 0);  -- csense_sdi:readdata -> mm_interconnect_2:csense_sdi_s1_readdata
	signal mm_interconnect_2_csense_sdi_s1_address                                                : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_sdi_s1_address -> csense_sdi:address
	signal mm_interconnect_2_csense_sdi_s1_write                                                  : std_logic;                      -- mm_interconnect_2:csense_sdi_s1_write -> mm_interconnect_2_csense_sdi_s1_write:in
	signal mm_interconnect_2_csense_sdi_s1_writedata                                              : std_logic_vector(31 downto 0);  -- mm_interconnect_2:csense_sdi_s1_writedata -> csense_sdi:writedata
	signal mm_interconnect_2_csense_sck_s1_chipselect                                             : std_logic;                      -- mm_interconnect_2:csense_sck_s1_chipselect -> csense_sck:chipselect
	signal mm_interconnect_2_csense_sck_s1_readdata                                               : std_logic_vector(31 downto 0);  -- csense_sck:readdata -> mm_interconnect_2:csense_sck_s1_readdata
	signal mm_interconnect_2_csense_sck_s1_address                                                : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_sck_s1_address -> csense_sck:address
	signal mm_interconnect_2_csense_sck_s1_write                                                  : std_logic;                      -- mm_interconnect_2:csense_sck_s1_write -> mm_interconnect_2_csense_sck_s1_write:in
	signal mm_interconnect_2_csense_sck_s1_writedata                                              : std_logic_vector(31 downto 0);  -- mm_interconnect_2:csense_sck_s1_writedata -> csense_sck:writedata
	signal mm_interconnect_2_csense_cs_n_s1_chipselect                                            : std_logic;                      -- mm_interconnect_2:csense_cs_n_s1_chipselect -> csense_cs_n:chipselect
	signal mm_interconnect_2_csense_cs_n_s1_readdata                                              : std_logic_vector(31 downto 0);  -- csense_cs_n:readdata -> mm_interconnect_2:csense_cs_n_s1_readdata
	signal mm_interconnect_2_csense_cs_n_s1_address                                               : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_cs_n_s1_address -> csense_cs_n:address
	signal mm_interconnect_2_csense_cs_n_s1_write                                                 : std_logic;                      -- mm_interconnect_2:csense_cs_n_s1_write -> mm_interconnect_2_csense_cs_n_s1_write:in
	signal mm_interconnect_2_csense_cs_n_s1_writedata                                             : std_logic_vector(31 downto 0);  -- mm_interconnect_2:csense_cs_n_s1_writedata -> csense_cs_n:writedata
	signal mm_interconnect_2_csense_adc_fo_s1_chipselect                                          : std_logic;                      -- mm_interconnect_2:csense_adc_fo_s1_chipselect -> csense_adc_fo:chipselect
	signal mm_interconnect_2_csense_adc_fo_s1_readdata                                            : std_logic_vector(31 downto 0);  -- csense_adc_fo:readdata -> mm_interconnect_2:csense_adc_fo_s1_readdata
	signal mm_interconnect_2_csense_adc_fo_s1_address                                             : std_logic_vector(1 downto 0);   -- mm_interconnect_2:csense_adc_fo_s1_address -> csense_adc_fo:address
	signal mm_interconnect_2_csense_adc_fo_s1_write                                               : std_logic;                      -- mm_interconnect_2:csense_adc_fo_s1_write -> mm_interconnect_2_csense_adc_fo_s1_write:in
	signal mm_interconnect_2_csense_adc_fo_s1_writedata                                           : std_logic_vector(31 downto 0);  -- mm_interconnect_2:csense_adc_fo_s1_writedata -> csense_adc_fo:writedata
	signal mm_interconnect_2_pio_led_painel_s1_chipselect                                         : std_logic;                      -- mm_interconnect_2:pio_LED_painel_s1_chipselect -> pio_LED_painel:chipselect
	signal mm_interconnect_2_pio_led_painel_s1_readdata                                           : std_logic_vector(31 downto 0);  -- pio_LED_painel:readdata -> mm_interconnect_2:pio_LED_painel_s1_readdata
	signal mm_interconnect_2_pio_led_painel_s1_address                                            : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_LED_painel_s1_address -> pio_LED_painel:address
	signal mm_interconnect_2_pio_led_painel_s1_write                                              : std_logic;                      -- mm_interconnect_2:pio_LED_painel_s1_write -> mm_interconnect_2_pio_led_painel_s1_write:in
	signal mm_interconnect_2_pio_led_painel_s1_writedata                                          : std_logic_vector(31 downto 0);  -- mm_interconnect_2:pio_LED_painel_s1_writedata -> pio_LED_painel:writedata
	signal mm_interconnect_2_rtcc_alarm_s1_readdata                                               : std_logic_vector(31 downto 0);  -- rtcc_alarm:readdata -> mm_interconnect_2:rtcc_alarm_s1_readdata
	signal mm_interconnect_2_rtcc_alarm_s1_address                                                : std_logic_vector(1 downto 0);   -- mm_interconnect_2:rtcc_alarm_s1_address -> rtcc_alarm:address
	signal mm_interconnect_2_rtcc_sdo_s1_readdata                                                 : std_logic_vector(31 downto 0);  -- rtcc_sdo:readdata -> mm_interconnect_2:rtcc_sdo_s1_readdata
	signal mm_interconnect_2_rtcc_sdo_s1_address                                                  : std_logic_vector(1 downto 0);   -- mm_interconnect_2:rtcc_sdo_s1_address -> rtcc_sdo:address
	signal mm_interconnect_2_rtcc_sdi_s1_chipselect                                               : std_logic;                      -- mm_interconnect_2:rtcc_sdi_s1_chipselect -> rtcc_sdi:chipselect
	signal mm_interconnect_2_rtcc_sdi_s1_readdata                                                 : std_logic_vector(31 downto 0);  -- rtcc_sdi:readdata -> mm_interconnect_2:rtcc_sdi_s1_readdata
	signal mm_interconnect_2_rtcc_sdi_s1_address                                                  : std_logic_vector(1 downto 0);   -- mm_interconnect_2:rtcc_sdi_s1_address -> rtcc_sdi:address
	signal mm_interconnect_2_rtcc_sdi_s1_write                                                    : std_logic;                      -- mm_interconnect_2:rtcc_sdi_s1_write -> mm_interconnect_2_rtcc_sdi_s1_write:in
	signal mm_interconnect_2_rtcc_sdi_s1_writedata                                                : std_logic_vector(31 downto 0);  -- mm_interconnect_2:rtcc_sdi_s1_writedata -> rtcc_sdi:writedata
	signal mm_interconnect_2_rtcc_sck_s1_chipselect                                               : std_logic;                      -- mm_interconnect_2:rtcc_sck_s1_chipselect -> rtcc_sck:chipselect
	signal mm_interconnect_2_rtcc_sck_s1_readdata                                                 : std_logic_vector(31 downto 0);  -- rtcc_sck:readdata -> mm_interconnect_2:rtcc_sck_s1_readdata
	signal mm_interconnect_2_rtcc_sck_s1_address                                                  : std_logic_vector(1 downto 0);   -- mm_interconnect_2:rtcc_sck_s1_address -> rtcc_sck:address
	signal mm_interconnect_2_rtcc_sck_s1_write                                                    : std_logic;                      -- mm_interconnect_2:rtcc_sck_s1_write -> mm_interconnect_2_rtcc_sck_s1_write:in
	signal mm_interconnect_2_rtcc_sck_s1_writedata                                                : std_logic_vector(31 downto 0);  -- mm_interconnect_2:rtcc_sck_s1_writedata -> rtcc_sck:writedata
	signal mm_interconnect_2_rtcc_cs_n_s1_chipselect                                              : std_logic;                      -- mm_interconnect_2:rtcc_cs_n_s1_chipselect -> rtcc_cs_n:chipselect
	signal mm_interconnect_2_rtcc_cs_n_s1_readdata                                                : std_logic_vector(31 downto 0);  -- rtcc_cs_n:readdata -> mm_interconnect_2:rtcc_cs_n_s1_readdata
	signal mm_interconnect_2_rtcc_cs_n_s1_address                                                 : std_logic_vector(1 downto 0);   -- mm_interconnect_2:rtcc_cs_n_s1_address -> rtcc_cs_n:address
	signal mm_interconnect_2_rtcc_cs_n_s1_write                                                   : std_logic;                      -- mm_interconnect_2:rtcc_cs_n_s1_write -> mm_interconnect_2_rtcc_cs_n_s1_write:in
	signal mm_interconnect_2_rtcc_cs_n_s1_writedata                                               : std_logic_vector(31 downto 0);  -- mm_interconnect_2:rtcc_cs_n_s1_writedata -> rtcc_cs_n:writedata
	signal mm_interconnect_2_rs232_uart_s1_chipselect                                             : std_logic;                      -- mm_interconnect_2:rs232_uart_s1_chipselect -> rs232_uart:chipselect
	signal mm_interconnect_2_rs232_uart_s1_readdata                                               : std_logic_vector(15 downto 0);  -- rs232_uart:readdata -> mm_interconnect_2:rs232_uart_s1_readdata
	signal mm_interconnect_2_rs232_uart_s1_address                                                : std_logic_vector(2 downto 0);   -- mm_interconnect_2:rs232_uart_s1_address -> rs232_uart:address
	signal mm_interconnect_2_rs232_uart_s1_read                                                   : std_logic;                      -- mm_interconnect_2:rs232_uart_s1_read -> mm_interconnect_2_rs232_uart_s1_read:in
	signal mm_interconnect_2_rs232_uart_s1_begintransfer                                          : std_logic;                      -- mm_interconnect_2:rs232_uart_s1_begintransfer -> rs232_uart:begintransfer
	signal mm_interconnect_2_rs232_uart_s1_write                                                  : std_logic;                      -- mm_interconnect_2:rs232_uart_s1_write -> mm_interconnect_2_rs232_uart_s1_write:in
	signal mm_interconnect_2_rs232_uart_s1_writedata                                              : std_logic_vector(15 downto 0);  -- mm_interconnect_2:rs232_uart_s1_writedata -> rs232_uart:writedata
	signal mm_interconnect_2_pio_ctrl_io_lvds_s1_chipselect                                       : std_logic;                      -- mm_interconnect_2:pio_ctrl_io_lvds_s1_chipselect -> pio_ctrl_io_lvds:chipselect
	signal mm_interconnect_2_pio_ctrl_io_lvds_s1_readdata                                         : std_logic_vector(31 downto 0);  -- pio_ctrl_io_lvds:readdata -> mm_interconnect_2:pio_ctrl_io_lvds_s1_readdata
	signal mm_interconnect_2_pio_ctrl_io_lvds_s1_address                                          : std_logic_vector(1 downto 0);   -- mm_interconnect_2:pio_ctrl_io_lvds_s1_address -> pio_ctrl_io_lvds:address
	signal mm_interconnect_2_pio_ctrl_io_lvds_s1_write                                            : std_logic;                      -- mm_interconnect_2:pio_ctrl_io_lvds_s1_write -> mm_interconnect_2_pio_ctrl_io_lvds_s1_write:in
	signal mm_interconnect_2_pio_ctrl_io_lvds_s1_writedata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_2:pio_ctrl_io_lvds_s1_writedata -> pio_ctrl_io_lvds:writedata
	signal m1_clock_bridge_m0_waitrequest                                                         : std_logic;                      -- mm_interconnect_3:m1_clock_bridge_m0_waitrequest -> m1_clock_bridge:m0_waitrequest
	signal m1_clock_bridge_m0_readdata                                                            : std_logic_vector(255 downto 0); -- mm_interconnect_3:m1_clock_bridge_m0_readdata -> m1_clock_bridge:m0_readdata
	signal m1_clock_bridge_m0_debugaccess                                                         : std_logic;                      -- m1_clock_bridge:m0_debugaccess -> mm_interconnect_3:m1_clock_bridge_m0_debugaccess
	signal m1_clock_bridge_m0_address                                                             : std_logic_vector(30 downto 0);  -- m1_clock_bridge:m0_address -> mm_interconnect_3:m1_clock_bridge_m0_address
	signal m1_clock_bridge_m0_read                                                                : std_logic;                      -- m1_clock_bridge:m0_read -> mm_interconnect_3:m1_clock_bridge_m0_read
	signal m1_clock_bridge_m0_byteenable                                                          : std_logic_vector(31 downto 0);  -- m1_clock_bridge:m0_byteenable -> mm_interconnect_3:m1_clock_bridge_m0_byteenable
	signal m1_clock_bridge_m0_readdatavalid                                                       : std_logic;                      -- mm_interconnect_3:m1_clock_bridge_m0_readdatavalid -> m1_clock_bridge:m0_readdatavalid
	signal m1_clock_bridge_m0_writedata                                                           : std_logic_vector(255 downto 0); -- m1_clock_bridge:m0_writedata -> mm_interconnect_3:m1_clock_bridge_m0_writedata
	signal m1_clock_bridge_m0_write                                                               : std_logic;                      -- m1_clock_bridge:m0_write -> mm_interconnect_3:m1_clock_bridge_m0_write
	signal m1_clock_bridge_m0_burstcount                                                          : std_logic_vector(2 downto 0);   -- m1_clock_bridge:m0_burstcount -> mm_interconnect_3:m1_clock_bridge_m0_burstcount
	signal mm_interconnect_3_m1_ddr2_memory_avl_beginbursttransfer                                : std_logic;                      -- mm_interconnect_3:m1_ddr2_memory_avl_beginbursttransfer -> m1_ddr2_memory:avl_burstbegin
	signal mm_interconnect_3_m1_ddr2_memory_avl_readdata                                          : std_logic_vector(255 downto 0); -- m1_ddr2_memory:avl_rdata -> mm_interconnect_3:m1_ddr2_memory_avl_readdata
	signal m1_ddr2_memory_avl_waitrequest                                                         : std_logic;                      -- m1_ddr2_memory:avl_ready -> m1_ddr2_memory_avl_waitrequest:in
	signal mm_interconnect_3_m1_ddr2_memory_avl_address                                           : std_logic_vector(25 downto 0);  -- mm_interconnect_3:m1_ddr2_memory_avl_address -> m1_ddr2_memory:avl_addr
	signal mm_interconnect_3_m1_ddr2_memory_avl_read                                              : std_logic;                      -- mm_interconnect_3:m1_ddr2_memory_avl_read -> m1_ddr2_memory:avl_read_req
	signal mm_interconnect_3_m1_ddr2_memory_avl_byteenable                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_3:m1_ddr2_memory_avl_byteenable -> m1_ddr2_memory:avl_be
	signal mm_interconnect_3_m1_ddr2_memory_avl_readdatavalid                                     : std_logic;                      -- m1_ddr2_memory:avl_rdata_valid -> mm_interconnect_3:m1_ddr2_memory_avl_readdatavalid
	signal mm_interconnect_3_m1_ddr2_memory_avl_write                                             : std_logic;                      -- mm_interconnect_3:m1_ddr2_memory_avl_write -> m1_ddr2_memory:avl_write_req
	signal mm_interconnect_3_m1_ddr2_memory_avl_writedata                                         : std_logic_vector(255 downto 0); -- mm_interconnect_3:m1_ddr2_memory_avl_writedata -> m1_ddr2_memory:avl_wdata
	signal mm_interconnect_3_m1_ddr2_memory_avl_burstcount                                        : std_logic_vector(7 downto 0);   -- mm_interconnect_3:m1_ddr2_memory_avl_burstcount -> m1_ddr2_memory:avl_size
	signal m1_ddr2_memory_afi_clk_clk                                                             : std_logic;                      -- m1_ddr2_memory:afi_clk -> [mm_interconnect_3:m1_ddr2_memory_afi_clk_clk, rst_controller_016:clk]
	signal dma_ftdi_usb3_mm_read_readdata                                                         : std_logic_vector(255 downto 0); -- mm_interconnect_4:dma_ftdi_usb3_mm_read_readdata -> dma_ftdi_usb3:mm_read_readdata
	signal dma_ftdi_usb3_mm_read_waitrequest                                                      : std_logic;                      -- mm_interconnect_4:dma_ftdi_usb3_mm_read_waitrequest -> dma_ftdi_usb3:mm_read_waitrequest
	signal dma_ftdi_usb3_mm_read_address                                                          : std_logic_vector(33 downto 0);  -- dma_ftdi_usb3:mm_read_address -> mm_interconnect_4:dma_ftdi_usb3_mm_read_address
	signal dma_ftdi_usb3_mm_read_read                                                             : std_logic;                      -- dma_ftdi_usb3:mm_read_read -> mm_interconnect_4:dma_ftdi_usb3_mm_read_read
	signal dma_ftdi_usb3_mm_read_byteenable                                                       : std_logic_vector(31 downto 0);  -- dma_ftdi_usb3:mm_read_byteenable -> mm_interconnect_4:dma_ftdi_usb3_mm_read_byteenable
	signal dma_ftdi_usb3_mm_read_readdatavalid                                                    : std_logic;                      -- mm_interconnect_4:dma_ftdi_usb3_mm_read_readdatavalid -> dma_ftdi_usb3:mm_read_readdatavalid
	signal mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_readdata                               : std_logic_vector(255 downto 0); -- FTDI_USB3_0:avalon_slave_data_readdata -> mm_interconnect_4:FTDI_USB3_0_avalon_slave_data_readdata
	signal mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_waitrequest                            : std_logic;                      -- FTDI_USB3_0:avalon_slave_data_waitrequest -> mm_interconnect_4:FTDI_USB3_0_avalon_slave_data_waitrequest
	signal mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_address                                : std_logic_vector(20 downto 0);  -- mm_interconnect_4:FTDI_USB3_0_avalon_slave_data_address -> FTDI_USB3_0:avalon_slave_data_address
	signal mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_read                                   : std_logic;                      -- mm_interconnect_4:FTDI_USB3_0_avalon_slave_data_read -> FTDI_USB3_0:avalon_slave_data_read
	signal mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_write                                  : std_logic;                      -- mm_interconnect_4:FTDI_USB3_0_avalon_slave_data_write -> FTDI_USB3_0:avalon_slave_data_write
	signal mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_writedata                              : std_logic_vector(255 downto 0); -- mm_interconnect_4:FTDI_USB3_0_avalon_slave_data_writedata -> FTDI_USB3_0:avalon_slave_data_writedata
	signal dma_comm_1_left_mm_write_waitrequest                                                   : std_logic;                      -- mm_interconnect_5:dma_comm_1_left_mm_write_waitrequest -> dma_comm_1_left:mm_write_waitrequest
	signal dma_comm_1_left_mm_write_address                                                       : std_logic_vector(32 downto 0);  -- dma_comm_1_left:mm_write_address -> mm_interconnect_5:dma_comm_1_left_mm_write_address
	signal dma_comm_1_left_mm_write_byteenable                                                    : std_logic_vector(31 downto 0);  -- dma_comm_1_left:mm_write_byteenable -> mm_interconnect_5:dma_comm_1_left_mm_write_byteenable
	signal dma_comm_1_left_mm_write_write                                                         : std_logic;                      -- dma_comm_1_left:mm_write_write -> mm_interconnect_5:dma_comm_1_left_mm_write_write
	signal dma_comm_1_left_mm_write_writedata                                                     : std_logic_vector(255 downto 0); -- dma_comm_1_left:mm_write_writedata -> mm_interconnect_5:dma_comm_1_left_mm_write_writedata
	signal mm_interconnect_5_comm_pedreiro_v1_01_a_avalon_slave_l_buffer_waitrequest              : std_logic;                      -- COMM_Pedreiro_v1_01_A:avalon_slave_L_buffer_waitrequest -> mm_interconnect_5:COMM_Pedreiro_v1_01_A_avalon_slave_L_buffer_waitrequest
	signal mm_interconnect_5_comm_pedreiro_v1_01_a_avalon_slave_l_buffer_address                  : std_logic_vector(20 downto 0);  -- mm_interconnect_5:COMM_Pedreiro_v1_01_A_avalon_slave_L_buffer_address -> COMM_Pedreiro_v1_01_A:avalon_slave_L_buffer_address
	signal mm_interconnect_5_comm_pedreiro_v1_01_a_avalon_slave_l_buffer_write                    : std_logic;                      -- mm_interconnect_5:COMM_Pedreiro_v1_01_A_avalon_slave_L_buffer_write -> COMM_Pedreiro_v1_01_A:avalon_slave_L_buffer_write
	signal mm_interconnect_5_comm_pedreiro_v1_01_a_avalon_slave_l_buffer_writedata                : std_logic_vector(255 downto 0); -- mm_interconnect_5:COMM_Pedreiro_v1_01_A_avalon_slave_L_buffer_writedata -> COMM_Pedreiro_v1_01_A:avalon_slave_L_buffer_writedata
	signal dma_comm_2_left_mm_write_waitrequest                                                   : std_logic;                      -- mm_interconnect_6:dma_comm_2_left_mm_write_waitrequest -> dma_comm_2_left:mm_write_waitrequest
	signal dma_comm_2_left_mm_write_address                                                       : std_logic_vector(32 downto 0);  -- dma_comm_2_left:mm_write_address -> mm_interconnect_6:dma_comm_2_left_mm_write_address
	signal dma_comm_2_left_mm_write_byteenable                                                    : std_logic_vector(31 downto 0);  -- dma_comm_2_left:mm_write_byteenable -> mm_interconnect_6:dma_comm_2_left_mm_write_byteenable
	signal dma_comm_2_left_mm_write_write                                                         : std_logic;                      -- dma_comm_2_left:mm_write_write -> mm_interconnect_6:dma_comm_2_left_mm_write_write
	signal dma_comm_2_left_mm_write_writedata                                                     : std_logic_vector(255 downto 0); -- dma_comm_2_left:mm_write_writedata -> mm_interconnect_6:dma_comm_2_left_mm_write_writedata
	signal mm_interconnect_6_comm_pedreiro_v1_01_b_avalon_slave_l_buffer_waitrequest              : std_logic;                      -- COMM_Pedreiro_v1_01_B:avalon_slave_L_buffer_waitrequest -> mm_interconnect_6:COMM_Pedreiro_v1_01_B_avalon_slave_L_buffer_waitrequest
	signal mm_interconnect_6_comm_pedreiro_v1_01_b_avalon_slave_l_buffer_address                  : std_logic_vector(20 downto 0);  -- mm_interconnect_6:COMM_Pedreiro_v1_01_B_avalon_slave_L_buffer_address -> COMM_Pedreiro_v1_01_B:avalon_slave_L_buffer_address
	signal mm_interconnect_6_comm_pedreiro_v1_01_b_avalon_slave_l_buffer_write                    : std_logic;                      -- mm_interconnect_6:COMM_Pedreiro_v1_01_B_avalon_slave_L_buffer_write -> COMM_Pedreiro_v1_01_B:avalon_slave_L_buffer_write
	signal mm_interconnect_6_comm_pedreiro_v1_01_b_avalon_slave_l_buffer_writedata                : std_logic_vector(255 downto 0); -- mm_interconnect_6:COMM_Pedreiro_v1_01_B_avalon_slave_L_buffer_writedata -> COMM_Pedreiro_v1_01_B:avalon_slave_L_buffer_writedata
	signal dma_comm_3_left_mm_write_waitrequest                                                   : std_logic;                      -- mm_interconnect_7:dma_comm_3_left_mm_write_waitrequest -> dma_comm_3_left:mm_write_waitrequest
	signal dma_comm_3_left_mm_write_address                                                       : std_logic_vector(32 downto 0);  -- dma_comm_3_left:mm_write_address -> mm_interconnect_7:dma_comm_3_left_mm_write_address
	signal dma_comm_3_left_mm_write_byteenable                                                    : std_logic_vector(31 downto 0);  -- dma_comm_3_left:mm_write_byteenable -> mm_interconnect_7:dma_comm_3_left_mm_write_byteenable
	signal dma_comm_3_left_mm_write_write                                                         : std_logic;                      -- dma_comm_3_left:mm_write_write -> mm_interconnect_7:dma_comm_3_left_mm_write_write
	signal dma_comm_3_left_mm_write_writedata                                                     : std_logic_vector(255 downto 0); -- dma_comm_3_left:mm_write_writedata -> mm_interconnect_7:dma_comm_3_left_mm_write_writedata
	signal mm_interconnect_7_comm_pedreiro_v1_01_c_avalon_slave_l_buffer_waitrequest              : std_logic;                      -- COMM_Pedreiro_v1_01_C:avalon_slave_L_buffer_waitrequest -> mm_interconnect_7:COMM_Pedreiro_v1_01_C_avalon_slave_L_buffer_waitrequest
	signal mm_interconnect_7_comm_pedreiro_v1_01_c_avalon_slave_l_buffer_address                  : std_logic_vector(20 downto 0);  -- mm_interconnect_7:COMM_Pedreiro_v1_01_C_avalon_slave_L_buffer_address -> COMM_Pedreiro_v1_01_C:avalon_slave_L_buffer_address
	signal mm_interconnect_7_comm_pedreiro_v1_01_c_avalon_slave_l_buffer_write                    : std_logic;                      -- mm_interconnect_7:COMM_Pedreiro_v1_01_C_avalon_slave_L_buffer_write -> COMM_Pedreiro_v1_01_C:avalon_slave_L_buffer_write
	signal mm_interconnect_7_comm_pedreiro_v1_01_c_avalon_slave_l_buffer_writedata                : std_logic_vector(255 downto 0); -- mm_interconnect_7:COMM_Pedreiro_v1_01_C_avalon_slave_L_buffer_writedata -> COMM_Pedreiro_v1_01_C:avalon_slave_L_buffer_writedata
	signal dma_comm_4_left_mm_write_waitrequest                                                   : std_logic;                      -- mm_interconnect_8:dma_comm_4_left_mm_write_waitrequest -> dma_comm_4_left:mm_write_waitrequest
	signal dma_comm_4_left_mm_write_address                                                       : std_logic_vector(32 downto 0);  -- dma_comm_4_left:mm_write_address -> mm_interconnect_8:dma_comm_4_left_mm_write_address
	signal dma_comm_4_left_mm_write_byteenable                                                    : std_logic_vector(31 downto 0);  -- dma_comm_4_left:mm_write_byteenable -> mm_interconnect_8:dma_comm_4_left_mm_write_byteenable
	signal dma_comm_4_left_mm_write_write                                                         : std_logic;                      -- dma_comm_4_left:mm_write_write -> mm_interconnect_8:dma_comm_4_left_mm_write_write
	signal dma_comm_4_left_mm_write_writedata                                                     : std_logic_vector(255 downto 0); -- dma_comm_4_left:mm_write_writedata -> mm_interconnect_8:dma_comm_4_left_mm_write_writedata
	signal mm_interconnect_8_comm_pedreiro_v1_01_d_avalon_slave_l_buffer_waitrequest              : std_logic;                      -- COMM_Pedreiro_v1_01_D:avalon_slave_L_buffer_waitrequest -> mm_interconnect_8:COMM_Pedreiro_v1_01_D_avalon_slave_L_buffer_waitrequest
	signal mm_interconnect_8_comm_pedreiro_v1_01_d_avalon_slave_l_buffer_address                  : std_logic_vector(20 downto 0);  -- mm_interconnect_8:COMM_Pedreiro_v1_01_D_avalon_slave_L_buffer_address -> COMM_Pedreiro_v1_01_D:avalon_slave_L_buffer_address
	signal mm_interconnect_8_comm_pedreiro_v1_01_d_avalon_slave_l_buffer_write                    : std_logic;                      -- mm_interconnect_8:COMM_Pedreiro_v1_01_D_avalon_slave_L_buffer_write -> COMM_Pedreiro_v1_01_D:avalon_slave_L_buffer_write
	signal mm_interconnect_8_comm_pedreiro_v1_01_d_avalon_slave_l_buffer_writedata                : std_logic_vector(255 downto 0); -- mm_interconnect_8:COMM_Pedreiro_v1_01_D_avalon_slave_L_buffer_writedata -> COMM_Pedreiro_v1_01_D:avalon_slave_L_buffer_writedata
	signal dma_comm_5_left_mm_write_waitrequest                                                   : std_logic;                      -- mm_interconnect_9:dma_comm_5_left_mm_write_waitrequest -> dma_comm_5_left:mm_write_waitrequest
	signal dma_comm_5_left_mm_write_address                                                       : std_logic_vector(32 downto 0);  -- dma_comm_5_left:mm_write_address -> mm_interconnect_9:dma_comm_5_left_mm_write_address
	signal dma_comm_5_left_mm_write_byteenable                                                    : std_logic_vector(31 downto 0);  -- dma_comm_5_left:mm_write_byteenable -> mm_interconnect_9:dma_comm_5_left_mm_write_byteenable
	signal dma_comm_5_left_mm_write_write                                                         : std_logic;                      -- dma_comm_5_left:mm_write_write -> mm_interconnect_9:dma_comm_5_left_mm_write_write
	signal dma_comm_5_left_mm_write_writedata                                                     : std_logic_vector(255 downto 0); -- dma_comm_5_left:mm_write_writedata -> mm_interconnect_9:dma_comm_5_left_mm_write_writedata
	signal mm_interconnect_9_comm_pedreiro_v1_01_e_avalon_slave_l_buffer_waitrequest              : std_logic;                      -- COMM_Pedreiro_v1_01_E:avalon_slave_L_buffer_waitrequest -> mm_interconnect_9:COMM_Pedreiro_v1_01_E_avalon_slave_L_buffer_waitrequest
	signal mm_interconnect_9_comm_pedreiro_v1_01_e_avalon_slave_l_buffer_address                  : std_logic_vector(20 downto 0);  -- mm_interconnect_9:COMM_Pedreiro_v1_01_E_avalon_slave_L_buffer_address -> COMM_Pedreiro_v1_01_E:avalon_slave_L_buffer_address
	signal mm_interconnect_9_comm_pedreiro_v1_01_e_avalon_slave_l_buffer_write                    : std_logic;                      -- mm_interconnect_9:COMM_Pedreiro_v1_01_E_avalon_slave_L_buffer_write -> COMM_Pedreiro_v1_01_E:avalon_slave_L_buffer_write
	signal mm_interconnect_9_comm_pedreiro_v1_01_e_avalon_slave_l_buffer_writedata                : std_logic_vector(255 downto 0); -- mm_interconnect_9:COMM_Pedreiro_v1_01_E_avalon_slave_L_buffer_writedata -> COMM_Pedreiro_v1_01_E:avalon_slave_L_buffer_writedata
	signal dma_comm_6_left_mm_write_waitrequest                                                   : std_logic;                      -- mm_interconnect_10:dma_comm_6_left_mm_write_waitrequest -> dma_comm_6_left:mm_write_waitrequest
	signal dma_comm_6_left_mm_write_address                                                       : std_logic_vector(32 downto 0);  -- dma_comm_6_left:mm_write_address -> mm_interconnect_10:dma_comm_6_left_mm_write_address
	signal dma_comm_6_left_mm_write_byteenable                                                    : std_logic_vector(31 downto 0);  -- dma_comm_6_left:mm_write_byteenable -> mm_interconnect_10:dma_comm_6_left_mm_write_byteenable
	signal dma_comm_6_left_mm_write_write                                                         : std_logic;                      -- dma_comm_6_left:mm_write_write -> mm_interconnect_10:dma_comm_6_left_mm_write_write
	signal dma_comm_6_left_mm_write_writedata                                                     : std_logic_vector(255 downto 0); -- dma_comm_6_left:mm_write_writedata -> mm_interconnect_10:dma_comm_6_left_mm_write_writedata
	signal mm_interconnect_10_comm_pedreiro_v1_01_f_avalon_slave_l_buffer_waitrequest             : std_logic;                      -- COMM_Pedreiro_v1_01_F:avalon_slave_L_buffer_waitrequest -> mm_interconnect_10:COMM_Pedreiro_v1_01_F_avalon_slave_L_buffer_waitrequest
	signal mm_interconnect_10_comm_pedreiro_v1_01_f_avalon_slave_l_buffer_address                 : std_logic_vector(20 downto 0);  -- mm_interconnect_10:COMM_Pedreiro_v1_01_F_avalon_slave_L_buffer_address -> COMM_Pedreiro_v1_01_F:avalon_slave_L_buffer_address
	signal mm_interconnect_10_comm_pedreiro_v1_01_f_avalon_slave_l_buffer_write                   : std_logic;                      -- mm_interconnect_10:COMM_Pedreiro_v1_01_F_avalon_slave_L_buffer_write -> COMM_Pedreiro_v1_01_F:avalon_slave_L_buffer_write
	signal mm_interconnect_10_comm_pedreiro_v1_01_f_avalon_slave_l_buffer_writedata               : std_logic_vector(255 downto 0); -- mm_interconnect_10:COMM_Pedreiro_v1_01_F_avalon_slave_L_buffer_writedata -> COMM_Pedreiro_v1_01_F:avalon_slave_L_buffer_writedata
	signal dma_comm_1_right_mm_write_waitrequest                                                  : std_logic;                      -- mm_interconnect_11:dma_comm_1_right_mm_write_waitrequest -> dma_comm_1_right:mm_write_waitrequest
	signal dma_comm_1_right_mm_write_address                                                      : std_logic_vector(32 downto 0);  -- dma_comm_1_right:mm_write_address -> mm_interconnect_11:dma_comm_1_right_mm_write_address
	signal dma_comm_1_right_mm_write_byteenable                                                   : std_logic_vector(31 downto 0);  -- dma_comm_1_right:mm_write_byteenable -> mm_interconnect_11:dma_comm_1_right_mm_write_byteenable
	signal dma_comm_1_right_mm_write_write                                                        : std_logic;                      -- dma_comm_1_right:mm_write_write -> mm_interconnect_11:dma_comm_1_right_mm_write_write
	signal dma_comm_1_right_mm_write_writedata                                                    : std_logic_vector(255 downto 0); -- dma_comm_1_right:mm_write_writedata -> mm_interconnect_11:dma_comm_1_right_mm_write_writedata
	signal mm_interconnect_11_comm_pedreiro_v1_01_a_avalon_slave_r_buffer_waitrequest             : std_logic;                      -- COMM_Pedreiro_v1_01_A:avalon_slave_R_buffer_waitrequest -> mm_interconnect_11:COMM_Pedreiro_v1_01_A_avalon_slave_R_buffer_waitrequest
	signal mm_interconnect_11_comm_pedreiro_v1_01_a_avalon_slave_r_buffer_address                 : std_logic_vector(20 downto 0);  -- mm_interconnect_11:COMM_Pedreiro_v1_01_A_avalon_slave_R_buffer_address -> COMM_Pedreiro_v1_01_A:avalon_slave_R_buffer_address
	signal mm_interconnect_11_comm_pedreiro_v1_01_a_avalon_slave_r_buffer_write                   : std_logic;                      -- mm_interconnect_11:COMM_Pedreiro_v1_01_A_avalon_slave_R_buffer_write -> COMM_Pedreiro_v1_01_A:avalon_slave_R_buffer_write
	signal mm_interconnect_11_comm_pedreiro_v1_01_a_avalon_slave_r_buffer_writedata               : std_logic_vector(255 downto 0); -- mm_interconnect_11:COMM_Pedreiro_v1_01_A_avalon_slave_R_buffer_writedata -> COMM_Pedreiro_v1_01_A:avalon_slave_R_buffer_writedata
	signal dma_comm_2_right_mm_write_waitrequest                                                  : std_logic;                      -- mm_interconnect_12:dma_comm_2_right_mm_write_waitrequest -> dma_comm_2_right:mm_write_waitrequest
	signal dma_comm_2_right_mm_write_address                                                      : std_logic_vector(32 downto 0);  -- dma_comm_2_right:mm_write_address -> mm_interconnect_12:dma_comm_2_right_mm_write_address
	signal dma_comm_2_right_mm_write_byteenable                                                   : std_logic_vector(31 downto 0);  -- dma_comm_2_right:mm_write_byteenable -> mm_interconnect_12:dma_comm_2_right_mm_write_byteenable
	signal dma_comm_2_right_mm_write_write                                                        : std_logic;                      -- dma_comm_2_right:mm_write_write -> mm_interconnect_12:dma_comm_2_right_mm_write_write
	signal dma_comm_2_right_mm_write_writedata                                                    : std_logic_vector(255 downto 0); -- dma_comm_2_right:mm_write_writedata -> mm_interconnect_12:dma_comm_2_right_mm_write_writedata
	signal mm_interconnect_12_comm_pedreiro_v1_01_b_avalon_slave_r_buffer_waitrequest             : std_logic;                      -- COMM_Pedreiro_v1_01_B:avalon_slave_R_buffer_waitrequest -> mm_interconnect_12:COMM_Pedreiro_v1_01_B_avalon_slave_R_buffer_waitrequest
	signal mm_interconnect_12_comm_pedreiro_v1_01_b_avalon_slave_r_buffer_address                 : std_logic_vector(20 downto 0);  -- mm_interconnect_12:COMM_Pedreiro_v1_01_B_avalon_slave_R_buffer_address -> COMM_Pedreiro_v1_01_B:avalon_slave_R_buffer_address
	signal mm_interconnect_12_comm_pedreiro_v1_01_b_avalon_slave_r_buffer_write                   : std_logic;                      -- mm_interconnect_12:COMM_Pedreiro_v1_01_B_avalon_slave_R_buffer_write -> COMM_Pedreiro_v1_01_B:avalon_slave_R_buffer_write
	signal mm_interconnect_12_comm_pedreiro_v1_01_b_avalon_slave_r_buffer_writedata               : std_logic_vector(255 downto 0); -- mm_interconnect_12:COMM_Pedreiro_v1_01_B_avalon_slave_R_buffer_writedata -> COMM_Pedreiro_v1_01_B:avalon_slave_R_buffer_writedata
	signal dma_comm_3_right_mm_write_waitrequest                                                  : std_logic;                      -- mm_interconnect_13:dma_comm_3_right_mm_write_waitrequest -> dma_comm_3_right:mm_write_waitrequest
	signal dma_comm_3_right_mm_write_address                                                      : std_logic_vector(32 downto 0);  -- dma_comm_3_right:mm_write_address -> mm_interconnect_13:dma_comm_3_right_mm_write_address
	signal dma_comm_3_right_mm_write_byteenable                                                   : std_logic_vector(31 downto 0);  -- dma_comm_3_right:mm_write_byteenable -> mm_interconnect_13:dma_comm_3_right_mm_write_byteenable
	signal dma_comm_3_right_mm_write_write                                                        : std_logic;                      -- dma_comm_3_right:mm_write_write -> mm_interconnect_13:dma_comm_3_right_mm_write_write
	signal dma_comm_3_right_mm_write_writedata                                                    : std_logic_vector(255 downto 0); -- dma_comm_3_right:mm_write_writedata -> mm_interconnect_13:dma_comm_3_right_mm_write_writedata
	signal mm_interconnect_13_comm_pedreiro_v1_01_c_avalon_slave_r_buffer_waitrequest             : std_logic;                      -- COMM_Pedreiro_v1_01_C:avalon_slave_R_buffer_waitrequest -> mm_interconnect_13:COMM_Pedreiro_v1_01_C_avalon_slave_R_buffer_waitrequest
	signal mm_interconnect_13_comm_pedreiro_v1_01_c_avalon_slave_r_buffer_address                 : std_logic_vector(20 downto 0);  -- mm_interconnect_13:COMM_Pedreiro_v1_01_C_avalon_slave_R_buffer_address -> COMM_Pedreiro_v1_01_C:avalon_slave_R_buffer_address
	signal mm_interconnect_13_comm_pedreiro_v1_01_c_avalon_slave_r_buffer_write                   : std_logic;                      -- mm_interconnect_13:COMM_Pedreiro_v1_01_C_avalon_slave_R_buffer_write -> COMM_Pedreiro_v1_01_C:avalon_slave_R_buffer_write
	signal mm_interconnect_13_comm_pedreiro_v1_01_c_avalon_slave_r_buffer_writedata               : std_logic_vector(255 downto 0); -- mm_interconnect_13:COMM_Pedreiro_v1_01_C_avalon_slave_R_buffer_writedata -> COMM_Pedreiro_v1_01_C:avalon_slave_R_buffer_writedata
	signal dma_comm_4_right_mm_write_waitrequest                                                  : std_logic;                      -- mm_interconnect_14:dma_comm_4_right_mm_write_waitrequest -> dma_comm_4_right:mm_write_waitrequest
	signal dma_comm_4_right_mm_write_address                                                      : std_logic_vector(32 downto 0);  -- dma_comm_4_right:mm_write_address -> mm_interconnect_14:dma_comm_4_right_mm_write_address
	signal dma_comm_4_right_mm_write_byteenable                                                   : std_logic_vector(31 downto 0);  -- dma_comm_4_right:mm_write_byteenable -> mm_interconnect_14:dma_comm_4_right_mm_write_byteenable
	signal dma_comm_4_right_mm_write_write                                                        : std_logic;                      -- dma_comm_4_right:mm_write_write -> mm_interconnect_14:dma_comm_4_right_mm_write_write
	signal dma_comm_4_right_mm_write_writedata                                                    : std_logic_vector(255 downto 0); -- dma_comm_4_right:mm_write_writedata -> mm_interconnect_14:dma_comm_4_right_mm_write_writedata
	signal mm_interconnect_14_comm_pedreiro_v1_01_d_avalon_slave_r_buffer_waitrequest             : std_logic;                      -- COMM_Pedreiro_v1_01_D:avalon_slave_R_buffer_waitrequest -> mm_interconnect_14:COMM_Pedreiro_v1_01_D_avalon_slave_R_buffer_waitrequest
	signal mm_interconnect_14_comm_pedreiro_v1_01_d_avalon_slave_r_buffer_address                 : std_logic_vector(20 downto 0);  -- mm_interconnect_14:COMM_Pedreiro_v1_01_D_avalon_slave_R_buffer_address -> COMM_Pedreiro_v1_01_D:avalon_slave_R_buffer_address
	signal mm_interconnect_14_comm_pedreiro_v1_01_d_avalon_slave_r_buffer_write                   : std_logic;                      -- mm_interconnect_14:COMM_Pedreiro_v1_01_D_avalon_slave_R_buffer_write -> COMM_Pedreiro_v1_01_D:avalon_slave_R_buffer_write
	signal mm_interconnect_14_comm_pedreiro_v1_01_d_avalon_slave_r_buffer_writedata               : std_logic_vector(255 downto 0); -- mm_interconnect_14:COMM_Pedreiro_v1_01_D_avalon_slave_R_buffer_writedata -> COMM_Pedreiro_v1_01_D:avalon_slave_R_buffer_writedata
	signal dma_comm_5_right_mm_write_waitrequest                                                  : std_logic;                      -- mm_interconnect_15:dma_comm_5_right_mm_write_waitrequest -> dma_comm_5_right:mm_write_waitrequest
	signal dma_comm_5_right_mm_write_address                                                      : std_logic_vector(32 downto 0);  -- dma_comm_5_right:mm_write_address -> mm_interconnect_15:dma_comm_5_right_mm_write_address
	signal dma_comm_5_right_mm_write_byteenable                                                   : std_logic_vector(31 downto 0);  -- dma_comm_5_right:mm_write_byteenable -> mm_interconnect_15:dma_comm_5_right_mm_write_byteenable
	signal dma_comm_5_right_mm_write_write                                                        : std_logic;                      -- dma_comm_5_right:mm_write_write -> mm_interconnect_15:dma_comm_5_right_mm_write_write
	signal dma_comm_5_right_mm_write_writedata                                                    : std_logic_vector(255 downto 0); -- dma_comm_5_right:mm_write_writedata -> mm_interconnect_15:dma_comm_5_right_mm_write_writedata
	signal mm_interconnect_15_comm_pedreiro_v1_01_e_avalon_slave_r_buffer_waitrequest             : std_logic;                      -- COMM_Pedreiro_v1_01_E:avalon_slave_R_buffer_waitrequest -> mm_interconnect_15:COMM_Pedreiro_v1_01_E_avalon_slave_R_buffer_waitrequest
	signal mm_interconnect_15_comm_pedreiro_v1_01_e_avalon_slave_r_buffer_address                 : std_logic_vector(20 downto 0);  -- mm_interconnect_15:COMM_Pedreiro_v1_01_E_avalon_slave_R_buffer_address -> COMM_Pedreiro_v1_01_E:avalon_slave_R_buffer_address
	signal mm_interconnect_15_comm_pedreiro_v1_01_e_avalon_slave_r_buffer_write                   : std_logic;                      -- mm_interconnect_15:COMM_Pedreiro_v1_01_E_avalon_slave_R_buffer_write -> COMM_Pedreiro_v1_01_E:avalon_slave_R_buffer_write
	signal mm_interconnect_15_comm_pedreiro_v1_01_e_avalon_slave_r_buffer_writedata               : std_logic_vector(255 downto 0); -- mm_interconnect_15:COMM_Pedreiro_v1_01_E_avalon_slave_R_buffer_writedata -> COMM_Pedreiro_v1_01_E:avalon_slave_R_buffer_writedata
	signal dma_comm_6_right_mm_write_waitrequest                                                  : std_logic;                      -- mm_interconnect_16:dma_comm_6_right_mm_write_waitrequest -> dma_comm_6_right:mm_write_waitrequest
	signal dma_comm_6_right_mm_write_address                                                      : std_logic_vector(32 downto 0);  -- dma_comm_6_right:mm_write_address -> mm_interconnect_16:dma_comm_6_right_mm_write_address
	signal dma_comm_6_right_mm_write_byteenable                                                   : std_logic_vector(31 downto 0);  -- dma_comm_6_right:mm_write_byteenable -> mm_interconnect_16:dma_comm_6_right_mm_write_byteenable
	signal dma_comm_6_right_mm_write_write                                                        : std_logic;                      -- dma_comm_6_right:mm_write_write -> mm_interconnect_16:dma_comm_6_right_mm_write_write
	signal dma_comm_6_right_mm_write_writedata                                                    : std_logic_vector(255 downto 0); -- dma_comm_6_right:mm_write_writedata -> mm_interconnect_16:dma_comm_6_right_mm_write_writedata
	signal mm_interconnect_16_comm_pedreiro_v1_01_f_avalon_slave_r_buffer_waitrequest             : std_logic;                      -- COMM_Pedreiro_v1_01_F:avalon_slave_R_buffer_waitrequest -> mm_interconnect_16:COMM_Pedreiro_v1_01_F_avalon_slave_R_buffer_waitrequest
	signal mm_interconnect_16_comm_pedreiro_v1_01_f_avalon_slave_r_buffer_address                 : std_logic_vector(20 downto 0);  -- mm_interconnect_16:COMM_Pedreiro_v1_01_F_avalon_slave_R_buffer_address -> COMM_Pedreiro_v1_01_F:avalon_slave_R_buffer_address
	signal mm_interconnect_16_comm_pedreiro_v1_01_f_avalon_slave_r_buffer_write                   : std_logic;                      -- mm_interconnect_16:COMM_Pedreiro_v1_01_F_avalon_slave_R_buffer_write -> COMM_Pedreiro_v1_01_F:avalon_slave_R_buffer_write
	signal mm_interconnect_16_comm_pedreiro_v1_01_f_avalon_slave_r_buffer_writedata               : std_logic_vector(255 downto 0); -- mm_interconnect_16:COMM_Pedreiro_v1_01_F_avalon_slave_R_buffer_writedata -> COMM_Pedreiro_v1_01_F:avalon_slave_R_buffer_writedata
	signal irq_mapper_receiver0_irq                                                               : std_logic;                      -- COMM_Pedreiro_v1_01_A:buffers_interrupt_sender_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                               : std_logic;                      -- COMM_Pedreiro_v1_01_B:buffers_interrupt_sender_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                               : std_logic;                      -- COMM_Pedreiro_v1_01_C:buffers_interrupt_sender_irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                               : std_logic;                      -- COMM_Pedreiro_v1_01_D:buffers_interrupt_sender_irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                                               : std_logic;                      -- COMM_Pedreiro_v1_01_E:buffers_interrupt_sender_irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                                               : std_logic;                      -- COMM_Pedreiro_v1_01_F:buffers_interrupt_sender_irq -> irq_mapper:receiver5_irq
	signal irq_mapper_receiver6_irq                                                               : std_logic;                      -- dma_comm_1_left:csr_irq_irq -> irq_mapper:receiver6_irq
	signal irq_mapper_receiver7_irq                                                               : std_logic;                      -- dma_comm_1_right:csr_irq_irq -> irq_mapper:receiver7_irq
	signal irq_mapper_receiver8_irq                                                               : std_logic;                      -- dma_comm_2_left:csr_irq_irq -> irq_mapper:receiver8_irq
	signal irq_mapper_receiver9_irq                                                               : std_logic;                      -- dma_comm_2_right:csr_irq_irq -> irq_mapper:receiver9_irq
	signal irq_mapper_receiver10_irq                                                              : std_logic;                      -- dma_comm_3_left:csr_irq_irq -> irq_mapper:receiver10_irq
	signal irq_mapper_receiver11_irq                                                              : std_logic;                      -- dma_comm_3_right:csr_irq_irq -> irq_mapper:receiver11_irq
	signal irq_mapper_receiver12_irq                                                              : std_logic;                      -- dma_comm_4_left:csr_irq_irq -> irq_mapper:receiver12_irq
	signal irq_mapper_receiver13_irq                                                              : std_logic;                      -- dma_comm_4_right:csr_irq_irq -> irq_mapper:receiver13_irq
	signal irq_mapper_receiver14_irq                                                              : std_logic;                      -- dma_comm_6_right:csr_irq_irq -> irq_mapper:receiver14_irq
	signal irq_mapper_receiver15_irq                                                              : std_logic;                      -- dma_comm_6_left:csr_irq_irq -> irq_mapper:receiver15_irq
	signal irq_mapper_receiver16_irq                                                              : std_logic;                      -- dma_comm_5_right:csr_irq_irq -> irq_mapper:receiver16_irq
	signal irq_mapper_receiver17_irq                                                              : std_logic;                      -- dma_comm_5_left:csr_irq_irq -> irq_mapper:receiver17_irq
	signal irq_mapper_receiver18_irq                                                              : std_logic;                      -- dma_ftdi_usb3:csr_irq_irq -> irq_mapper:receiver18_irq
	signal irq_mapper_receiver19_irq                                                              : std_logic;                      -- FTDI_USB3_0:ftdi_interrupt_sender_irq -> irq_mapper:receiver19_irq
	signal irq_mapper_receiver20_irq                                                              : std_logic;                      -- jtag_uart_0:av_irq -> irq_mapper:receiver20_irq
	signal irq_mapper_receiver25_irq                                                              : std_logic;                      -- COMM_Pedreiro_v1_01_A:rmap_interrupt_sender_irq -> irq_mapper:receiver25_irq
	signal irq_mapper_receiver26_irq                                                              : std_logic;                      -- COMM_Pedreiro_v1_01_B:rmap_interrupt_sender_irq -> irq_mapper:receiver26_irq
	signal irq_mapper_receiver27_irq                                                              : std_logic;                      -- COMM_Pedreiro_v1_01_C:rmap_interrupt_sender_irq -> irq_mapper:receiver27_irq
	signal irq_mapper_receiver28_irq                                                              : std_logic;                      -- COMM_Pedreiro_v1_01_D:rmap_interrupt_sender_irq -> irq_mapper:receiver28_irq
	signal irq_mapper_receiver29_irq                                                              : std_logic;                      -- COMM_Pedreiro_v1_01_E:rmap_interrupt_sender_irq -> irq_mapper:receiver29_irq
	signal irq_mapper_receiver30_irq                                                              : std_logic;                      -- COMM_Pedreiro_v1_01_F:rmap_interrupt_sender_irq -> irq_mapper:receiver30_irq
	signal nios2_gen2_0_irq_irq                                                                   : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal irq_mapper_receiver21_irq                                                              : std_logic;                      -- irq_synchronizer:sender_irq -> irq_mapper:receiver21_irq
	signal irq_synchronizer_receiver_irq                                                          : std_logic_vector(0 downto 0);   -- timer_1ms:irq -> irq_synchronizer:receiver_irq
	signal irq_mapper_receiver22_irq                                                              : std_logic;                      -- irq_synchronizer_001:sender_irq -> irq_mapper:receiver22_irq
	signal irq_synchronizer_001_receiver_irq                                                      : std_logic_vector(0 downto 0);   -- timer_1us:irq -> irq_synchronizer_001:receiver_irq
	signal irq_mapper_receiver23_irq                                                              : std_logic;                      -- irq_synchronizer_002:sender_irq -> irq_mapper:receiver23_irq
	signal irq_synchronizer_002_receiver_irq                                                      : std_logic_vector(0 downto 0);   -- rs232_uart:irq -> irq_synchronizer_002:receiver_irq
	signal irq_mapper_receiver24_irq                                                              : std_logic;                      -- irq_synchronizer_003:sender_irq -> irq_mapper:receiver24_irq
	signal irq_synchronizer_003_receiver_irq                                                      : std_logic_vector(0 downto 0);   -- sync:pre_sync_interrupt_sender_irq_o -> irq_synchronizer_003:receiver_irq
	signal irq_mapper_receiver31_irq                                                              : std_logic;                      -- irq_synchronizer_004:sender_irq -> irq_mapper:receiver31_irq
	signal irq_synchronizer_004_receiver_irq                                                      : std_logic_vector(0 downto 0);   -- sync:sync_interrupt_sender_irq_o -> irq_synchronizer_004:receiver_irq
	signal rst_controller_001_reset_out_reset                                                     : std_logic;                      -- rst_controller_001:reset_out -> [mm_interconnect_2:Altera_UP_SD_Card_Avalon_Interface_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_reset_source_sd_card_reset                                              : std_logic;                      -- rst_controller:reset_source_sd_card_reset -> rst_controller_001:reset_in1
	signal rst_controller_002_reset_out_reset                                                     : std_logic;                      -- rst_controller_002:reset_out -> [COMM_Pedreiro_v1_01_A:reset_sink_reset, mm_interconnect_0:rmap_mem_nfee_comm_1_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_11:COMM_Pedreiro_v1_01_A_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:rmap_mem_nfee_comm_1_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_5:COMM_Pedreiro_v1_01_A_reset_sink_reset_bridge_in_reset_reset, rmap_mem_nfee_comm_1:reset_i]
	signal rst_controller_reset_source_comm_ch1_reset                                             : std_logic;                      -- rst_controller:reset_source_comm_ch1_reset -> rst_controller_002:reset_in1
	signal rst_controller_003_reset_out_reset                                                     : std_logic;                      -- rst_controller_003:reset_out -> [COMM_Pedreiro_v1_01_B:reset_sink_reset, mm_interconnect_0:rmap_mem_nfee_comm_2_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_12:COMM_Pedreiro_v1_01_B_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:rmap_mem_nfee_comm_2_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_6:COMM_Pedreiro_v1_01_B_reset_sink_reset_bridge_in_reset_reset, rmap_mem_nfee_comm_2:reset_i]
	signal rst_controller_reset_source_comm_ch2_reset                                             : std_logic;                      -- rst_controller:reset_source_comm_ch2_reset -> rst_controller_003:reset_in1
	signal rst_controller_004_reset_out_reset                                                     : std_logic;                      -- rst_controller_004:reset_out -> [COMM_Pedreiro_v1_01_C:reset_sink_reset, mm_interconnect_0:rmap_mem_nfee_comm_3_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_13:COMM_Pedreiro_v1_01_C_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:rmap_mem_nfee_comm_3_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_7:COMM_Pedreiro_v1_01_C_reset_sink_reset_bridge_in_reset_reset, rmap_mem_nfee_comm_3:reset_i]
	signal rst_controller_reset_source_comm_ch3_reset                                             : std_logic;                      -- rst_controller:reset_source_comm_ch3_reset -> rst_controller_004:reset_in1
	signal rst_controller_005_reset_out_reset                                                     : std_logic;                      -- rst_controller_005:reset_out -> [COMM_Pedreiro_v1_01_D:reset_sink_reset, mm_interconnect_0:rmap_mem_nfee_comm_4_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_14:COMM_Pedreiro_v1_01_D_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:rmap_mem_nfee_comm_4_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_8:COMM_Pedreiro_v1_01_D_reset_sink_reset_bridge_in_reset_reset, rmap_mem_nfee_comm_4:reset_i]
	signal rst_controller_reset_source_comm_ch4_reset                                             : std_logic;                      -- rst_controller:reset_source_comm_ch4_reset -> rst_controller_005:reset_in1
	signal rst_controller_006_reset_out_reset                                                     : std_logic;                      -- rst_controller_006:reset_out -> [COMM_Pedreiro_v1_01_E:reset_sink_reset, mm_interconnect_0:rmap_mem_nfee_comm_5_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_15:COMM_Pedreiro_v1_01_E_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:rmap_mem_nfee_comm_5_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_9:COMM_Pedreiro_v1_01_E_reset_sink_reset_bridge_in_reset_reset, rmap_mem_nfee_comm_5:reset_i]
	signal rst_controller_reset_source_comm_ch5_reset                                             : std_logic;                      -- rst_controller:reset_source_comm_ch5_reset -> rst_controller_006:reset_in1
	signal rst_controller_007_reset_out_reset                                                     : std_logic;                      -- rst_controller_007:reset_out -> [COMM_Pedreiro_v1_01_F:reset_sink_reset, mm_interconnect_0:rmap_mem_nfee_comm_6_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_10:COMM_Pedreiro_v1_01_F_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_16:COMM_Pedreiro_v1_01_F_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:rmap_mem_nfee_comm_6_reset_sink_reset_bridge_in_reset_reset, rmap_mem_nfee_comm_6:reset_i]
	signal rst_controller_reset_source_comm_ch6_reset                                             : std_logic;                      -- rst_controller:reset_source_comm_ch6_reset -> rst_controller_007:reset_in1
	signal rst_controller_008_reset_out_reset                                                     : std_logic;                      -- rst_controller_008:reset_out -> [FTDI_USB3_0:reset_sink_reset, clock_bridge_afi_50:s0_reset, ddr2_address_span_extender:reset, m1_clock_bridge:s0_reset, mm_interconnect_0:ddr2_address_span_extender_reset_reset_bridge_in_reset_reset, mm_interconnect_0:m1_clock_bridge_s0_reset_reset_bridge_in_reset_reset, mm_interconnect_10:dma_comm_6_left_reset_n_reset_bridge_in_reset_reset, mm_interconnect_11:dma_comm_1_right_reset_n_reset_bridge_in_reset_reset, mm_interconnect_12:dma_comm_2_right_reset_n_reset_bridge_in_reset_reset, mm_interconnect_13:dma_comm_3_right_reset_n_reset_bridge_in_reset_reset, mm_interconnect_14:dma_comm_4_right_reset_n_reset_bridge_in_reset_reset, mm_interconnect_15:dma_comm_5_right_reset_n_reset_bridge_in_reset_reset, mm_interconnect_16:dma_comm_6_right_reset_n_reset_bridge_in_reset_reset, mm_interconnect_1:jtag_uart_0_reset_reset_bridge_in_reset_reset, mm_interconnect_4:dma_ftdi_usb3_reset_n_reset_bridge_in_reset_reset, mm_interconnect_5:dma_comm_1_left_reset_n_reset_bridge_in_reset_reset, mm_interconnect_6:dma_comm_2_left_reset_n_reset_bridge_in_reset_reset, mm_interconnect_7:dma_comm_3_left_reset_n_reset_bridge_in_reset_reset, mm_interconnect_8:dma_comm_4_left_reset_n_reset_bridge_in_reset_reset, mm_interconnect_9:dma_comm_5_left_reset_n_reset_bridge_in_reset_reset, onchip_memory:reset, rst_controller_008_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_008_reset_out_reset_req                                                 : std_logic;                      -- rst_controller_008:reset_req -> [onchip_memory:reset_req, rst_translator:reset_req_in]
	signal rst_controller_009_reset_out_reset                                                     : std_logic;                      -- rst_controller_009:reset_out -> [SEVEN_SEGMENT_CONTROLLER_0:RST, clock_bridge_afi_50:m0_reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, mm_interconnect_2:clock_bridge_afi_50_m0_reset_reset_bridge_in_reset_reset, rst_controller:reset_sink_reset, rst_controller_009_reset_out_reset:in]
	signal rst_controller_010_reset_out_reset                                                     : std_logic;                      -- rst_controller_010:reset_out -> [ext_flash:reset_reset, mm_interconnect_1:ext_flash_reset_reset_bridge_in_reset_reset, tristate_conduit_bridge_0:reset]
	signal rst_controller_011_reset_out_reset                                                     : std_logic;                      -- rst_controller_011:reset_out -> [m1_clock_bridge:m0_reset, mm_interconnect_3:m1_clock_bridge_m0_reset_reset_bridge_in_reset_reset]
	signal rst_controller_012_reset_out_reset                                                     : std_logic;                      -- rst_controller_012:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, mm_interconnect_1:nios2_gen2_0_reset_reset_bridge_in_reset_reset, rst_controller_012_reset_out_reset:in, rst_translator_001:in_reset]
	signal rst_controller_012_reset_out_reset_req                                                 : std_logic;                      -- rst_controller_012:reset_req -> [nios2_gen2_0:reset_req, rst_translator_001:reset_req_in]
	signal rst_controller_013_reset_out_reset                                                     : std_logic;                      -- rst_controller_013:reset_out -> [irq_synchronizer_002:receiver_reset, mm_interconnect_2:rs232_uart_reset_reset_bridge_in_reset_reset, rst_controller_013_reset_out_reset:in]
	signal rst_controller_reset_source_rs232_reset                                                : std_logic;                      -- rst_controller:reset_source_rs232_reset -> rst_controller_013:reset_in1
	signal rst_controller_014_reset_out_reset                                                     : std_logic;                      -- rst_controller_014:reset_out -> [irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, mm_interconnect_2:sync_reset_reset_bridge_in_reset_reset, sync:reset_sink_reset_i]
	signal rst_controller_reset_source_sync_reset                                                 : std_logic;                      -- rst_controller:reset_source_sync_reset -> rst_controller_014:reset_in1
	signal rst_controller_015_reset_out_reset                                                     : std_logic;                      -- rst_controller_015:reset_out -> [mm_interconnect_0:m2_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:m2_ddr2_memory_soft_reset_reset_bridge_in_reset_reset]
	signal rst_controller_016_reset_out_reset                                                     : std_logic;                      -- rst_controller_016:reset_out -> [mm_interconnect_3:m1_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_3:m1_ddr2_memory_soft_reset_reset_bridge_in_reset_reset]
	signal rst_reset_n_ports_inv                                                                  : std_logic;                      -- rst_reset_n:inv -> [rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0, rst_controller_005:reset_in0, rst_controller_006:reset_in0, rst_controller_007:reset_in0, rst_controller_008:reset_in0, rst_controller_009:reset_in0, rst_controller_010:reset_in0, rst_controller_010:reset_in1, rst_controller_011:reset_in0, rst_controller_012:reset_in0, rst_controller_013:reset_in0, rst_controller_014:reset_in0, rst_controller_015:reset_in0, rst_controller_016:reset_in0]
	signal mm_interconnect_0_m2_ddr2_memory_avl_inv                                               : std_logic;                      -- m2_ddr2_memory_avl_waitrequest:inv -> mm_interconnect_0:m2_ddr2_memory_avl_waitrequest
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv                         : std_logic;                      -- mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv                        : std_logic;                      -- mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_2_m1_ddr2_i2c_sda_s1_write_ports_inv                                   : std_logic;                      -- mm_interconnect_2_m1_ddr2_i2c_sda_s1_write:inv -> m1_ddr2_i2c_sda:write_n
	signal mm_interconnect_2_m1_ddr2_i2c_scl_s1_write_ports_inv                                   : std_logic;                      -- mm_interconnect_2_m1_ddr2_i2c_scl_s1_write:inv -> m1_ddr2_i2c_scl:write_n
	signal mm_interconnect_2_pio_led_s1_write_ports_inv                                           : std_logic;                      -- mm_interconnect_2_pio_led_s1_write:inv -> pio_LED:write_n
	signal mm_interconnect_2_timer_1ms_s1_write_ports_inv                                         : std_logic;                      -- mm_interconnect_2_timer_1ms_s1_write:inv -> timer_1ms:write_n
	signal mm_interconnect_2_timer_1us_s1_write_ports_inv                                         : std_logic;                      -- mm_interconnect_2_timer_1us_s1_write:inv -> timer_1us:write_n
	signal mm_interconnect_2_temp_scl_s1_write_ports_inv                                          : std_logic;                      -- mm_interconnect_2_temp_scl_s1_write:inv -> temp_scl:write_n
	signal mm_interconnect_2_temp_sda_s1_write_ports_inv                                          : std_logic;                      -- mm_interconnect_2_temp_sda_s1_write:inv -> temp_sda:write_n
	signal mm_interconnect_2_m2_ddr2_i2c_sda_s1_write_ports_inv                                   : std_logic;                      -- mm_interconnect_2_m2_ddr2_i2c_sda_s1_write:inv -> m2_ddr2_i2c_sda:write_n
	signal mm_interconnect_2_m2_ddr2_i2c_scl_s1_write_ports_inv                                   : std_logic;                      -- mm_interconnect_2_m2_ddr2_i2c_scl_s1_write:inv -> m2_ddr2_i2c_scl:write_n
	signal mm_interconnect_2_csense_sdi_s1_write_ports_inv                                        : std_logic;                      -- mm_interconnect_2_csense_sdi_s1_write:inv -> csense_sdi:write_n
	signal mm_interconnect_2_csense_sck_s1_write_ports_inv                                        : std_logic;                      -- mm_interconnect_2_csense_sck_s1_write:inv -> csense_sck:write_n
	signal mm_interconnect_2_csense_cs_n_s1_write_ports_inv                                       : std_logic;                      -- mm_interconnect_2_csense_cs_n_s1_write:inv -> csense_cs_n:write_n
	signal mm_interconnect_2_csense_adc_fo_s1_write_ports_inv                                     : std_logic;                      -- mm_interconnect_2_csense_adc_fo_s1_write:inv -> csense_adc_fo:write_n
	signal mm_interconnect_2_pio_led_painel_s1_write_ports_inv                                    : std_logic;                      -- mm_interconnect_2_pio_led_painel_s1_write:inv -> pio_LED_painel:write_n
	signal mm_interconnect_2_rtcc_sdi_s1_write_ports_inv                                          : std_logic;                      -- mm_interconnect_2_rtcc_sdi_s1_write:inv -> rtcc_sdi:write_n
	signal mm_interconnect_2_rtcc_sck_s1_write_ports_inv                                          : std_logic;                      -- mm_interconnect_2_rtcc_sck_s1_write:inv -> rtcc_sck:write_n
	signal mm_interconnect_2_rtcc_cs_n_s1_write_ports_inv                                         : std_logic;                      -- mm_interconnect_2_rtcc_cs_n_s1_write:inv -> rtcc_cs_n:write_n
	signal mm_interconnect_2_rs232_uart_s1_read_ports_inv                                         : std_logic;                      -- mm_interconnect_2_rs232_uart_s1_read:inv -> rs232_uart:read_n
	signal mm_interconnect_2_rs232_uart_s1_write_ports_inv                                        : std_logic;                      -- mm_interconnect_2_rs232_uart_s1_write:inv -> rs232_uart:write_n
	signal mm_interconnect_2_pio_ctrl_io_lvds_s1_write_ports_inv                                  : std_logic;                      -- mm_interconnect_2_pio_ctrl_io_lvds_s1_write:inv -> pio_ctrl_io_lvds:write_n
	signal mm_interconnect_3_m1_ddr2_memory_avl_inv                                               : std_logic;                      -- m1_ddr2_memory_avl_waitrequest:inv -> mm_interconnect_3:m1_ddr2_memory_avl_waitrequest
	signal rst_controller_001_reset_out_reset_ports_inv                                           : std_logic;                      -- rst_controller_001_reset_out_reset:inv -> Altera_UP_SD_Card_Avalon_Interface_0:i_reset_n
	signal rst_controller_008_reset_out_reset_ports_inv                                           : std_logic;                      -- rst_controller_008_reset_out_reset:inv -> [dma_comm_1_left:reset_n_reset_n, dma_comm_1_right:reset_n_reset_n, dma_comm_2_left:reset_n_reset_n, dma_comm_2_right:reset_n_reset_n, dma_comm_3_left:reset_n_reset_n, dma_comm_3_right:reset_n_reset_n, dma_comm_4_left:reset_n_reset_n, dma_comm_4_right:reset_n_reset_n, dma_comm_5_left:reset_n_reset_n, dma_comm_5_right:reset_n_reset_n, dma_comm_6_left:reset_n_reset_n, dma_comm_6_right:reset_n_reset_n, dma_ftdi_usb3:reset_n_reset_n, jtag_uart_0:rst_n, sysid_qsys:reset_n]
	signal rst_controller_009_reset_out_reset_ports_inv                                           : std_logic;                      -- rst_controller_009_reset_out_reset:inv -> [csense_adc_fo:reset_n, csense_cs_n:reset_n, csense_sck:reset_n, csense_sdi:reset_n, csense_sdo:reset_n, m1_ddr2_i2c_scl:reset_n, m1_ddr2_i2c_sda:reset_n, m2_ddr2_i2c_scl:reset_n, m2_ddr2_i2c_sda:reset_n, pio_BUTTON:reset_n, pio_DIP:reset_n, pio_EXT:reset_n, pio_LED:reset_n, pio_LED_painel:reset_n, pio_ctrl_io_lvds:reset_n, rtcc_alarm:reset_n, rtcc_cs_n:reset_n, rtcc_sck:reset_n, rtcc_sdi:reset_n, rtcc_sdo:reset_n, sd_card_wp_n:reset_n, temp_scl:reset_n, temp_sda:reset_n, timer_1ms:reset_n, timer_1us:reset_n]
	signal rst_controller_012_reset_out_reset_ports_inv                                           : std_logic;                      -- rst_controller_012_reset_out_reset:inv -> nios2_gen2_0:reset_n
	signal rst_controller_013_reset_out_reset_ports_inv                                           : std_logic;                      -- rst_controller_013_reset_out_reset:inv -> rs232_uart:reset_n

begin

	altera_up_sd_card_avalon_interface_0 : component Altera_UP_SD_Card_Avalon_Interface
		port map (
			i_avalon_chip_select => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect,  -- avalon_sdcard_slave.chipselect
			i_avalon_address     => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address,     --                    .address
			i_avalon_read        => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read,        --                    .read
			i_avalon_write       => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write,       --                    .write
			i_avalon_byteenable  => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable,  --                    .byteenable
			i_avalon_writedata   => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata,   --                    .writedata
			o_avalon_readdata    => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata,    --                    .readdata
			o_avalon_waitrequest => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest, --                    .waitrequest
			i_clock              => clk50_clk,                                                                              --                 clk.clk
			i_reset_n            => rst_controller_001_reset_out_reset_ports_inv,                                           --               reset.reset_n
			b_SD_cmd             => sd_card_ip_b_SD_cmd,                                                                    --         conduit_end.export
			b_SD_dat             => sd_card_ip_b_SD_dat,                                                                    --                    .export
			b_SD_dat3            => sd_card_ip_b_SD_dat3,                                                                   --                    .export
			o_SD_clock           => sd_card_ip_o_SD_clock                                                                   --                    .export
		);

	comm_pedreiro_v1_01_a : component comm_v1_80_top
		port map (
			reset_sink_reset                   => rst_controller_002_reset_out_reset,                                           --                        reset_sink.reset
			data_in                            => comm_a_conduit_end_data_in_signal,                                            --                   spw_conduit_end.data_in_signal
			data_out                           => comm_a_conduit_end_data_out_signal,                                           --                                  .data_out_signal
			strobe_in                          => comm_a_conduit_end_strobe_in_signal,                                          --                                  .strobe_in_signal
			strobe_out                         => comm_a_conduit_end_strobe_out_signal,                                         --                                  .strobe_out_signal
			sync_channel                       => comm_a_sync_end_sync_channel_signal,                                          --                  sync_conduit_end.sync_channel_signal
			rmap_interrupt_sender_irq          => irq_mapper_receiver25_irq,                                                    --             rmap_interrupt_sender.irq
			buffers_interrupt_sender_irq       => irq_mapper_receiver0_irq,                                                     --          buffers_interrupt_sender.irq
			clock_sink_100_clk                 => m2_ddr2_memory_afi_half_clk_clk,                                              --                    clock_sink_100.clk
			clock_sink_200_clk                 => m2_ddr2_memory_afi_clk_clk,                                                   --                    clock_sink_200.clk
			avalon_slave_windowing_address     => mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_address,       --            avalon_slave_windowing.address
			avalon_slave_windowing_write       => mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_write,         --                                  .write
			avalon_slave_windowing_read        => mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_read,          --                                  .read
			avalon_slave_windowing_writedata   => mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_writedata,     --                                  .writedata
			avalon_slave_windowing_byteenable  => mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_byteenable,    --                                  .byteenable
			avalon_slave_windowing_readdata    => mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_readdata,      --                                  .readdata
			avalon_slave_windowing_waitrequest => mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_waitrequest,   --                                  .waitrequest
			avalon_slave_L_buffer_address      => mm_interconnect_5_comm_pedreiro_v1_01_a_avalon_slave_l_buffer_address,        --             avalon_slave_L_buffer.address
			avalon_slave_L_buffer_waitrequest  => mm_interconnect_5_comm_pedreiro_v1_01_a_avalon_slave_l_buffer_waitrequest,    --                                  .waitrequest
			avalon_slave_L_buffer_write        => mm_interconnect_5_comm_pedreiro_v1_01_a_avalon_slave_l_buffer_write,          --                                  .write
			avalon_slave_L_buffer_writedata    => mm_interconnect_5_comm_pedreiro_v1_01_a_avalon_slave_l_buffer_writedata,      --                                  .writedata
			avalon_slave_R_buffer_address      => mm_interconnect_11_comm_pedreiro_v1_01_a_avalon_slave_r_buffer_address,       --             avalon_slave_R_buffer.address
			avalon_slave_R_buffer_write        => mm_interconnect_11_comm_pedreiro_v1_01_a_avalon_slave_r_buffer_write,         --                                  .write
			avalon_slave_R_buffer_writedata    => mm_interconnect_11_comm_pedreiro_v1_01_a_avalon_slave_r_buffer_writedata,     --                                  .writedata
			avalon_slave_R_buffer_waitrequest  => mm_interconnect_11_comm_pedreiro_v1_01_a_avalon_slave_r_buffer_waitrequest,   --                                  .waitrequest
			measurements_channel               => comm_a_measurements_conduit_end_measurements_channel_signal,                  --          measurements_conduit_end.measurements_channel_signal
			fee_codec_rmap_wr_waitrequest_i    => rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal,      -- conduit_end_fee_rmap_master_codec.wr_waitrequest_signal
			fee_codec_rmap_readdata_i          => rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_readdata_signal,            --                                  .readdata_signal
			fee_codec_rmap_rd_waitrequest_i    => rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal,      --                                  .rd_waitrequest_signal
			fee_codec_rmap_wr_address_o        => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_wr_address_signal,    --                                  .wr_address_signal
			fee_codec_rmap_write_o             => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_write_signal,         --                                  .write_signal
			fee_codec_rmap_writedata_o         => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_writedata_signal,     --                                  .writedata_signal
			fee_codec_rmap_rd_address_o        => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_rd_address_signal,    --                                  .rd_address_signal
			fee_codec_rmap_read_o              => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_read_signal,          --                                  .read_signal
			fee_hk_rmap_wr_waitrequest_i       => rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal,      --    conduit_end_fee_rmap_master_hk.wr_waitrequest_signal
			fee_hk_rmap_readdata_i             => rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_readdata_signal,            --                                  .readdata_signal
			fee_hk_rmap_rd_waitrequest_i       => rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal,      --                                  .rd_waitrequest_signal
			fee_hk_rmap_wr_address_o           => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_wr_address_signal,       --                                  .wr_address_signal
			fee_hk_rmap_write_o                => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_write_signal,            --                                  .write_signal
			fee_hk_rmap_writedata_o            => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_writedata_signal,        --                                  .writedata_signal
			fee_hk_rmap_rd_address_o           => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_rd_address_signal,       --                                  .rd_address_signal
			fee_hk_rmap_read_o                 => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_read_signal,             --                                  .read_signal
			channel_hk_timecode_control_o      => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_timecode_control_signal,     --        conduit_end_channel_hk_out.timecode_control_signal
			channel_hk_timecode_time_o         => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_timecode_time_signal,        --                                  .timecode_time_signal
			channel_hk_rmap_target_status_o    => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_rmap_target_status_signal,   --                                  .rmap_target_status_signal
			channel_hk_rmap_target_indicate_o  => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_rmap_target_indicate_signal, --                                  .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_o   => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_escape_err_signal,  --                                  .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_o   => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_credit_err_signal,  --                                  .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_o   => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_parity_err_signal,  --                                  .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_o   => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_disconnect_signal,  --                                  .spw_link_disconnect_signal
			channel_hk_spw_link_running_o      => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_running_signal,     --                                  .spw_link_running_signal
			channel_hk_frame_counter_o         => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_frame_counter_signal,        --                                  .frame_counter_signal
			channel_hk_frame_number_o          => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_frame_number_signal,         --                                  .frame_number_signal
			channel_win_mem_addr_offset_o      => comm_pedreiro_v1_01_a_conduit_end_avm_configs_out_win_mem_addr_offset_signal  --       conduit_end_avm_configs_out.win_mem_addr_offset_signal
		);

	comm_pedreiro_v1_01_b : component comm_v1_80_top
		port map (
			reset_sink_reset                   => rst_controller_003_reset_out_reset,                                           --                        reset_sink.reset
			data_in                            => comm_b_conduit_end_data_in_signal,                                            --                   spw_conduit_end.data_in_signal
			data_out                           => comm_b_conduit_end_data_out_signal,                                           --                                  .data_out_signal
			strobe_in                          => comm_b_conduit_end_strobe_in_signal,                                          --                                  .strobe_in_signal
			strobe_out                         => comm_b_conduit_end_strobe_out_signal,                                         --                                  .strobe_out_signal
			sync_channel                       => comm_b_sync_end_sync_channel_signal,                                          --                  sync_conduit_end.sync_channel_signal
			rmap_interrupt_sender_irq          => irq_mapper_receiver26_irq,                                                    --             rmap_interrupt_sender.irq
			buffers_interrupt_sender_irq       => irq_mapper_receiver1_irq,                                                     --          buffers_interrupt_sender.irq
			clock_sink_100_clk                 => m2_ddr2_memory_afi_half_clk_clk,                                              --                    clock_sink_100.clk
			clock_sink_200_clk                 => m2_ddr2_memory_afi_clk_clk,                                                   --                    clock_sink_200.clk
			avalon_slave_windowing_address     => mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_address,       --            avalon_slave_windowing.address
			avalon_slave_windowing_write       => mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_write,         --                                  .write
			avalon_slave_windowing_read        => mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_read,          --                                  .read
			avalon_slave_windowing_writedata   => mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_writedata,     --                                  .writedata
			avalon_slave_windowing_byteenable  => mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_byteenable,    --                                  .byteenable
			avalon_slave_windowing_readdata    => mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_readdata,      --                                  .readdata
			avalon_slave_windowing_waitrequest => mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_waitrequest,   --                                  .waitrequest
			avalon_slave_L_buffer_address      => mm_interconnect_6_comm_pedreiro_v1_01_b_avalon_slave_l_buffer_address,        --             avalon_slave_L_buffer.address
			avalon_slave_L_buffer_waitrequest  => mm_interconnect_6_comm_pedreiro_v1_01_b_avalon_slave_l_buffer_waitrequest,    --                                  .waitrequest
			avalon_slave_L_buffer_write        => mm_interconnect_6_comm_pedreiro_v1_01_b_avalon_slave_l_buffer_write,          --                                  .write
			avalon_slave_L_buffer_writedata    => mm_interconnect_6_comm_pedreiro_v1_01_b_avalon_slave_l_buffer_writedata,      --                                  .writedata
			avalon_slave_R_buffer_address      => mm_interconnect_12_comm_pedreiro_v1_01_b_avalon_slave_r_buffer_address,       --             avalon_slave_R_buffer.address
			avalon_slave_R_buffer_write        => mm_interconnect_12_comm_pedreiro_v1_01_b_avalon_slave_r_buffer_write,         --                                  .write
			avalon_slave_R_buffer_writedata    => mm_interconnect_12_comm_pedreiro_v1_01_b_avalon_slave_r_buffer_writedata,     --                                  .writedata
			avalon_slave_R_buffer_waitrequest  => mm_interconnect_12_comm_pedreiro_v1_01_b_avalon_slave_r_buffer_waitrequest,   --                                  .waitrequest
			measurements_channel               => comm_b_measurements_conduit_end_measurements_channel_signal,                  --          measurements_conduit_end.measurements_channel_signal
			fee_codec_rmap_wr_waitrequest_i    => rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal,      -- conduit_end_fee_rmap_master_codec.wr_waitrequest_signal
			fee_codec_rmap_readdata_i          => rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_readdata_signal,            --                                  .readdata_signal
			fee_codec_rmap_rd_waitrequest_i    => rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal,      --                                  .rd_waitrequest_signal
			fee_codec_rmap_wr_address_o        => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_wr_address_signal,    --                                  .wr_address_signal
			fee_codec_rmap_write_o             => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_write_signal,         --                                  .write_signal
			fee_codec_rmap_writedata_o         => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_writedata_signal,     --                                  .writedata_signal
			fee_codec_rmap_rd_address_o        => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_rd_address_signal,    --                                  .rd_address_signal
			fee_codec_rmap_read_o              => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_read_signal,          --                                  .read_signal
			fee_hk_rmap_wr_waitrequest_i       => rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal,      --    conduit_end_fee_rmap_master_hk.wr_waitrequest_signal
			fee_hk_rmap_readdata_i             => rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_readdata_signal,            --                                  .readdata_signal
			fee_hk_rmap_rd_waitrequest_i       => rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal,      --                                  .rd_waitrequest_signal
			fee_hk_rmap_wr_address_o           => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_wr_address_signal,       --                                  .wr_address_signal
			fee_hk_rmap_write_o                => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_write_signal,            --                                  .write_signal
			fee_hk_rmap_writedata_o            => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_writedata_signal,        --                                  .writedata_signal
			fee_hk_rmap_rd_address_o           => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_rd_address_signal,       --                                  .rd_address_signal
			fee_hk_rmap_read_o                 => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_read_signal,             --                                  .read_signal
			channel_hk_timecode_control_o      => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_timecode_control_signal,     --        conduit_end_channel_hk_out.timecode_control_signal
			channel_hk_timecode_time_o         => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_timecode_time_signal,        --                                  .timecode_time_signal
			channel_hk_rmap_target_status_o    => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_rmap_target_status_signal,   --                                  .rmap_target_status_signal
			channel_hk_rmap_target_indicate_o  => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_rmap_target_indicate_signal, --                                  .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_o   => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_escape_err_signal,  --                                  .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_o   => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_credit_err_signal,  --                                  .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_o   => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_parity_err_signal,  --                                  .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_o   => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_disconnect_signal,  --                                  .spw_link_disconnect_signal
			channel_hk_spw_link_running_o      => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_running_signal,     --                                  .spw_link_running_signal
			channel_hk_frame_counter_o         => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_frame_counter_signal,        --                                  .frame_counter_signal
			channel_hk_frame_number_o          => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_frame_number_signal,         --                                  .frame_number_signal
			channel_win_mem_addr_offset_o      => comm_pedreiro_v1_01_b_conduit_end_avm_configs_out_win_mem_addr_offset_signal  --       conduit_end_avm_configs_out.win_mem_addr_offset_signal
		);

	comm_pedreiro_v1_01_c : component comm_v1_80_top
		port map (
			reset_sink_reset                   => rst_controller_004_reset_out_reset,                                           --                        reset_sink.reset
			data_in                            => comm_c_conduit_end_data_in_signal,                                            --                   spw_conduit_end.data_in_signal
			data_out                           => comm_c_conduit_end_data_out_signal,                                           --                                  .data_out_signal
			strobe_in                          => comm_c_conduit_end_strobe_in_signal,                                          --                                  .strobe_in_signal
			strobe_out                         => comm_c_conduit_end_strobe_out_signal,                                         --                                  .strobe_out_signal
			sync_channel                       => comm_c_sync_end_sync_channel_signal,                                          --                  sync_conduit_end.sync_channel_signal
			rmap_interrupt_sender_irq          => irq_mapper_receiver27_irq,                                                    --             rmap_interrupt_sender.irq
			buffers_interrupt_sender_irq       => irq_mapper_receiver2_irq,                                                     --          buffers_interrupt_sender.irq
			clock_sink_100_clk                 => m2_ddr2_memory_afi_half_clk_clk,                                              --                    clock_sink_100.clk
			clock_sink_200_clk                 => m2_ddr2_memory_afi_clk_clk,                                                   --                    clock_sink_200.clk
			avalon_slave_windowing_address     => mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_address,       --            avalon_slave_windowing.address
			avalon_slave_windowing_write       => mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_write,         --                                  .write
			avalon_slave_windowing_read        => mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_read,          --                                  .read
			avalon_slave_windowing_writedata   => mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_writedata,     --                                  .writedata
			avalon_slave_windowing_byteenable  => mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_byteenable,    --                                  .byteenable
			avalon_slave_windowing_readdata    => mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_readdata,      --                                  .readdata
			avalon_slave_windowing_waitrequest => mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_waitrequest,   --                                  .waitrequest
			avalon_slave_L_buffer_address      => mm_interconnect_7_comm_pedreiro_v1_01_c_avalon_slave_l_buffer_address,        --             avalon_slave_L_buffer.address
			avalon_slave_L_buffer_waitrequest  => mm_interconnect_7_comm_pedreiro_v1_01_c_avalon_slave_l_buffer_waitrequest,    --                                  .waitrequest
			avalon_slave_L_buffer_write        => mm_interconnect_7_comm_pedreiro_v1_01_c_avalon_slave_l_buffer_write,          --                                  .write
			avalon_slave_L_buffer_writedata    => mm_interconnect_7_comm_pedreiro_v1_01_c_avalon_slave_l_buffer_writedata,      --                                  .writedata
			avalon_slave_R_buffer_address      => mm_interconnect_13_comm_pedreiro_v1_01_c_avalon_slave_r_buffer_address,       --             avalon_slave_R_buffer.address
			avalon_slave_R_buffer_write        => mm_interconnect_13_comm_pedreiro_v1_01_c_avalon_slave_r_buffer_write,         --                                  .write
			avalon_slave_R_buffer_writedata    => mm_interconnect_13_comm_pedreiro_v1_01_c_avalon_slave_r_buffer_writedata,     --                                  .writedata
			avalon_slave_R_buffer_waitrequest  => mm_interconnect_13_comm_pedreiro_v1_01_c_avalon_slave_r_buffer_waitrequest,   --                                  .waitrequest
			measurements_channel               => comm_c_measurements_conduit_end_measurements_channel_signal,                  --          measurements_conduit_end.measurements_channel_signal
			fee_codec_rmap_wr_waitrequest_i    => rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal,      -- conduit_end_fee_rmap_master_codec.wr_waitrequest_signal
			fee_codec_rmap_readdata_i          => rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_readdata_signal,            --                                  .readdata_signal
			fee_codec_rmap_rd_waitrequest_i    => rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal,      --                                  .rd_waitrequest_signal
			fee_codec_rmap_wr_address_o        => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_wr_address_signal,    --                                  .wr_address_signal
			fee_codec_rmap_write_o             => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_write_signal,         --                                  .write_signal
			fee_codec_rmap_writedata_o         => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_writedata_signal,     --                                  .writedata_signal
			fee_codec_rmap_rd_address_o        => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_rd_address_signal,    --                                  .rd_address_signal
			fee_codec_rmap_read_o              => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_read_signal,          --                                  .read_signal
			fee_hk_rmap_wr_waitrequest_i       => rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal,      --    conduit_end_fee_rmap_master_hk.wr_waitrequest_signal
			fee_hk_rmap_readdata_i             => rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_readdata_signal,            --                                  .readdata_signal
			fee_hk_rmap_rd_waitrequest_i       => rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal,      --                                  .rd_waitrequest_signal
			fee_hk_rmap_wr_address_o           => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_wr_address_signal,       --                                  .wr_address_signal
			fee_hk_rmap_write_o                => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_write_signal,            --                                  .write_signal
			fee_hk_rmap_writedata_o            => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_writedata_signal,        --                                  .writedata_signal
			fee_hk_rmap_rd_address_o           => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_rd_address_signal,       --                                  .rd_address_signal
			fee_hk_rmap_read_o                 => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_read_signal,             --                                  .read_signal
			channel_hk_timecode_control_o      => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_timecode_control_signal,     --        conduit_end_channel_hk_out.timecode_control_signal
			channel_hk_timecode_time_o         => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_timecode_time_signal,        --                                  .timecode_time_signal
			channel_hk_rmap_target_status_o    => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_rmap_target_status_signal,   --                                  .rmap_target_status_signal
			channel_hk_rmap_target_indicate_o  => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_rmap_target_indicate_signal, --                                  .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_o   => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_escape_err_signal,  --                                  .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_o   => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_credit_err_signal,  --                                  .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_o   => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_parity_err_signal,  --                                  .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_o   => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_disconnect_signal,  --                                  .spw_link_disconnect_signal
			channel_hk_spw_link_running_o      => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_running_signal,     --                                  .spw_link_running_signal
			channel_hk_frame_counter_o         => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_frame_counter_signal,        --                                  .frame_counter_signal
			channel_hk_frame_number_o          => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_frame_number_signal,         --                                  .frame_number_signal
			channel_win_mem_addr_offset_o      => comm_pedreiro_v1_01_c_conduit_end_avm_configs_out_win_mem_addr_offset_signal  --       conduit_end_avm_configs_out.win_mem_addr_offset_signal
		);

	comm_pedreiro_v1_01_d : component comm_v1_80_top
		port map (
			reset_sink_reset                   => rst_controller_005_reset_out_reset,                                           --                        reset_sink.reset
			data_in                            => comm_d_conduit_end_data_in_signal,                                            --                   spw_conduit_end.data_in_signal
			data_out                           => comm_d_conduit_end_data_out_signal,                                           --                                  .data_out_signal
			strobe_in                          => comm_d_conduit_end_strobe_in_signal,                                          --                                  .strobe_in_signal
			strobe_out                         => comm_d_conduit_end_strobe_out_signal,                                         --                                  .strobe_out_signal
			sync_channel                       => comm_d_sync_end_sync_channel_signal,                                          --                  sync_conduit_end.sync_channel_signal
			rmap_interrupt_sender_irq          => irq_mapper_receiver28_irq,                                                    --             rmap_interrupt_sender.irq
			buffers_interrupt_sender_irq       => irq_mapper_receiver3_irq,                                                     --          buffers_interrupt_sender.irq
			clock_sink_100_clk                 => m2_ddr2_memory_afi_half_clk_clk,                                              --                    clock_sink_100.clk
			clock_sink_200_clk                 => m2_ddr2_memory_afi_clk_clk,                                                   --                    clock_sink_200.clk
			avalon_slave_windowing_address     => mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_address,       --            avalon_slave_windowing.address
			avalon_slave_windowing_write       => mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_write,         --                                  .write
			avalon_slave_windowing_read        => mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_read,          --                                  .read
			avalon_slave_windowing_writedata   => mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_writedata,     --                                  .writedata
			avalon_slave_windowing_byteenable  => mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_byteenable,    --                                  .byteenable
			avalon_slave_windowing_readdata    => mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_readdata,      --                                  .readdata
			avalon_slave_windowing_waitrequest => mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_waitrequest,   --                                  .waitrequest
			avalon_slave_L_buffer_address      => mm_interconnect_8_comm_pedreiro_v1_01_d_avalon_slave_l_buffer_address,        --             avalon_slave_L_buffer.address
			avalon_slave_L_buffer_waitrequest  => mm_interconnect_8_comm_pedreiro_v1_01_d_avalon_slave_l_buffer_waitrequest,    --                                  .waitrequest
			avalon_slave_L_buffer_write        => mm_interconnect_8_comm_pedreiro_v1_01_d_avalon_slave_l_buffer_write,          --                                  .write
			avalon_slave_L_buffer_writedata    => mm_interconnect_8_comm_pedreiro_v1_01_d_avalon_slave_l_buffer_writedata,      --                                  .writedata
			avalon_slave_R_buffer_address      => mm_interconnect_14_comm_pedreiro_v1_01_d_avalon_slave_r_buffer_address,       --             avalon_slave_R_buffer.address
			avalon_slave_R_buffer_write        => mm_interconnect_14_comm_pedreiro_v1_01_d_avalon_slave_r_buffer_write,         --                                  .write
			avalon_slave_R_buffer_writedata    => mm_interconnect_14_comm_pedreiro_v1_01_d_avalon_slave_r_buffer_writedata,     --                                  .writedata
			avalon_slave_R_buffer_waitrequest  => mm_interconnect_14_comm_pedreiro_v1_01_d_avalon_slave_r_buffer_waitrequest,   --                                  .waitrequest
			measurements_channel               => comm_d_measurements_conduit_end_measurements_channel_signal,                  --          measurements_conduit_end.measurements_channel_signal
			fee_codec_rmap_wr_waitrequest_i    => rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal,      -- conduit_end_fee_rmap_master_codec.wr_waitrequest_signal
			fee_codec_rmap_readdata_i          => rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_readdata_signal,            --                                  .readdata_signal
			fee_codec_rmap_rd_waitrequest_i    => rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal,      --                                  .rd_waitrequest_signal
			fee_codec_rmap_wr_address_o        => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_wr_address_signal,    --                                  .wr_address_signal
			fee_codec_rmap_write_o             => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_write_signal,         --                                  .write_signal
			fee_codec_rmap_writedata_o         => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_writedata_signal,     --                                  .writedata_signal
			fee_codec_rmap_rd_address_o        => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_rd_address_signal,    --                                  .rd_address_signal
			fee_codec_rmap_read_o              => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_read_signal,          --                                  .read_signal
			fee_hk_rmap_wr_waitrequest_i       => rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal,      --    conduit_end_fee_rmap_master_hk.wr_waitrequest_signal
			fee_hk_rmap_readdata_i             => rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_readdata_signal,            --                                  .readdata_signal
			fee_hk_rmap_rd_waitrequest_i       => rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal,      --                                  .rd_waitrequest_signal
			fee_hk_rmap_wr_address_o           => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_wr_address_signal,       --                                  .wr_address_signal
			fee_hk_rmap_write_o                => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_write_signal,            --                                  .write_signal
			fee_hk_rmap_writedata_o            => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_writedata_signal,        --                                  .writedata_signal
			fee_hk_rmap_rd_address_o           => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_rd_address_signal,       --                                  .rd_address_signal
			fee_hk_rmap_read_o                 => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_read_signal,             --                                  .read_signal
			channel_hk_timecode_control_o      => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_timecode_control_signal,     --        conduit_end_channel_hk_out.timecode_control_signal
			channel_hk_timecode_time_o         => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_timecode_time_signal,        --                                  .timecode_time_signal
			channel_hk_rmap_target_status_o    => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_rmap_target_status_signal,   --                                  .rmap_target_status_signal
			channel_hk_rmap_target_indicate_o  => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_rmap_target_indicate_signal, --                                  .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_o   => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_escape_err_signal,  --                                  .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_o   => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_credit_err_signal,  --                                  .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_o   => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_parity_err_signal,  --                                  .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_o   => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_disconnect_signal,  --                                  .spw_link_disconnect_signal
			channel_hk_spw_link_running_o      => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_running_signal,     --                                  .spw_link_running_signal
			channel_hk_frame_counter_o         => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_frame_counter_signal,        --                                  .frame_counter_signal
			channel_hk_frame_number_o          => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_frame_number_signal,         --                                  .frame_number_signal
			channel_win_mem_addr_offset_o      => comm_pedreiro_v1_01_d_conduit_end_avm_configs_out_win_mem_addr_offset_signal  --       conduit_end_avm_configs_out.win_mem_addr_offset_signal
		);

	comm_pedreiro_v1_01_e : component comm_v1_80_top
		port map (
			reset_sink_reset                   => rst_controller_006_reset_out_reset,                                           --                        reset_sink.reset
			data_in                            => comm_e_conduit_end_data_in_signal,                                            --                   spw_conduit_end.data_in_signal
			data_out                           => comm_e_conduit_end_data_out_signal,                                           --                                  .data_out_signal
			strobe_in                          => comm_e_conduit_end_strobe_in_signal,                                          --                                  .strobe_in_signal
			strobe_out                         => comm_e_conduit_end_strobe_out_signal,                                         --                                  .strobe_out_signal
			sync_channel                       => comm_e_sync_end_sync_channel_signal,                                          --                  sync_conduit_end.sync_channel_signal
			rmap_interrupt_sender_irq          => irq_mapper_receiver29_irq,                                                    --             rmap_interrupt_sender.irq
			buffers_interrupt_sender_irq       => irq_mapper_receiver4_irq,                                                     --          buffers_interrupt_sender.irq
			clock_sink_100_clk                 => m2_ddr2_memory_afi_half_clk_clk,                                              --                    clock_sink_100.clk
			clock_sink_200_clk                 => m2_ddr2_memory_afi_clk_clk,                                                   --                    clock_sink_200.clk
			avalon_slave_windowing_address     => mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_address,       --            avalon_slave_windowing.address
			avalon_slave_windowing_write       => mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_write,         --                                  .write
			avalon_slave_windowing_read        => mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_read,          --                                  .read
			avalon_slave_windowing_writedata   => mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_writedata,     --                                  .writedata
			avalon_slave_windowing_byteenable  => mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_byteenable,    --                                  .byteenable
			avalon_slave_windowing_readdata    => mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_readdata,      --                                  .readdata
			avalon_slave_windowing_waitrequest => mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_waitrequest,   --                                  .waitrequest
			avalon_slave_L_buffer_address      => mm_interconnect_9_comm_pedreiro_v1_01_e_avalon_slave_l_buffer_address,        --             avalon_slave_L_buffer.address
			avalon_slave_L_buffer_waitrequest  => mm_interconnect_9_comm_pedreiro_v1_01_e_avalon_slave_l_buffer_waitrequest,    --                                  .waitrequest
			avalon_slave_L_buffer_write        => mm_interconnect_9_comm_pedreiro_v1_01_e_avalon_slave_l_buffer_write,          --                                  .write
			avalon_slave_L_buffer_writedata    => mm_interconnect_9_comm_pedreiro_v1_01_e_avalon_slave_l_buffer_writedata,      --                                  .writedata
			avalon_slave_R_buffer_address      => mm_interconnect_15_comm_pedreiro_v1_01_e_avalon_slave_r_buffer_address,       --             avalon_slave_R_buffer.address
			avalon_slave_R_buffer_write        => mm_interconnect_15_comm_pedreiro_v1_01_e_avalon_slave_r_buffer_write,         --                                  .write
			avalon_slave_R_buffer_writedata    => mm_interconnect_15_comm_pedreiro_v1_01_e_avalon_slave_r_buffer_writedata,     --                                  .writedata
			avalon_slave_R_buffer_waitrequest  => mm_interconnect_15_comm_pedreiro_v1_01_e_avalon_slave_r_buffer_waitrequest,   --                                  .waitrequest
			measurements_channel               => comm_e_measurements_conduit_end_measurements_channel_signal,                  --          measurements_conduit_end.measurements_channel_signal
			fee_codec_rmap_wr_waitrequest_i    => rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal,      -- conduit_end_fee_rmap_master_codec.wr_waitrequest_signal
			fee_codec_rmap_readdata_i          => rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_readdata_signal,            --                                  .readdata_signal
			fee_codec_rmap_rd_waitrequest_i    => rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal,      --                                  .rd_waitrequest_signal
			fee_codec_rmap_wr_address_o        => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_wr_address_signal,    --                                  .wr_address_signal
			fee_codec_rmap_write_o             => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_write_signal,         --                                  .write_signal
			fee_codec_rmap_writedata_o         => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_writedata_signal,     --                                  .writedata_signal
			fee_codec_rmap_rd_address_o        => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_rd_address_signal,    --                                  .rd_address_signal
			fee_codec_rmap_read_o              => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_read_signal,          --                                  .read_signal
			fee_hk_rmap_wr_waitrequest_i       => rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal,      --    conduit_end_fee_rmap_master_hk.wr_waitrequest_signal
			fee_hk_rmap_readdata_i             => rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_readdata_signal,            --                                  .readdata_signal
			fee_hk_rmap_rd_waitrequest_i       => rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal,      --                                  .rd_waitrequest_signal
			fee_hk_rmap_wr_address_o           => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_wr_address_signal,       --                                  .wr_address_signal
			fee_hk_rmap_write_o                => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_write_signal,            --                                  .write_signal
			fee_hk_rmap_writedata_o            => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_writedata_signal,        --                                  .writedata_signal
			fee_hk_rmap_rd_address_o           => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_rd_address_signal,       --                                  .rd_address_signal
			fee_hk_rmap_read_o                 => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_read_signal,             --                                  .read_signal
			channel_hk_timecode_control_o      => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_timecode_control_signal,     --        conduit_end_channel_hk_out.timecode_control_signal
			channel_hk_timecode_time_o         => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_timecode_time_signal,        --                                  .timecode_time_signal
			channel_hk_rmap_target_status_o    => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_rmap_target_status_signal,   --                                  .rmap_target_status_signal
			channel_hk_rmap_target_indicate_o  => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_rmap_target_indicate_signal, --                                  .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_o   => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_escape_err_signal,  --                                  .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_o   => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_credit_err_signal,  --                                  .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_o   => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_parity_err_signal,  --                                  .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_o   => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_disconnect_signal,  --                                  .spw_link_disconnect_signal
			channel_hk_spw_link_running_o      => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_running_signal,     --                                  .spw_link_running_signal
			channel_hk_frame_counter_o         => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_frame_counter_signal,        --                                  .frame_counter_signal
			channel_hk_frame_number_o          => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_frame_number_signal,         --                                  .frame_number_signal
			channel_win_mem_addr_offset_o      => comm_pedreiro_v1_01_e_conduit_end_avm_configs_out_win_mem_addr_offset_signal  --       conduit_end_avm_configs_out.win_mem_addr_offset_signal
		);

	comm_pedreiro_v1_01_f : component comm_v1_80_top
		port map (
			reset_sink_reset                   => rst_controller_007_reset_out_reset,                                           --                        reset_sink.reset
			data_in                            => comm_f_conduit_end_data_in_signal,                                            --                   spw_conduit_end.data_in_signal
			data_out                           => comm_f_conduit_end_data_out_signal,                                           --                                  .data_out_signal
			strobe_in                          => comm_f_conduit_end_strobe_in_signal,                                          --                                  .strobe_in_signal
			strobe_out                         => comm_f_conduit_end_strobe_out_signal,                                         --                                  .strobe_out_signal
			sync_channel                       => comm_f_sync_end_sync_channel_signal,                                          --                  sync_conduit_end.sync_channel_signal
			rmap_interrupt_sender_irq          => irq_mapper_receiver30_irq,                                                    --             rmap_interrupt_sender.irq
			buffers_interrupt_sender_irq       => irq_mapper_receiver5_irq,                                                     --          buffers_interrupt_sender.irq
			clock_sink_100_clk                 => m2_ddr2_memory_afi_half_clk_clk,                                              --                    clock_sink_100.clk
			clock_sink_200_clk                 => m2_ddr2_memory_afi_clk_clk,                                                   --                    clock_sink_200.clk
			avalon_slave_windowing_address     => mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_address,       --            avalon_slave_windowing.address
			avalon_slave_windowing_write       => mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_write,         --                                  .write
			avalon_slave_windowing_read        => mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_read,          --                                  .read
			avalon_slave_windowing_writedata   => mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_writedata,     --                                  .writedata
			avalon_slave_windowing_byteenable  => mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_byteenable,    --                                  .byteenable
			avalon_slave_windowing_readdata    => mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_readdata,      --                                  .readdata
			avalon_slave_windowing_waitrequest => mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_waitrequest,   --                                  .waitrequest
			avalon_slave_L_buffer_address      => mm_interconnect_10_comm_pedreiro_v1_01_f_avalon_slave_l_buffer_address,       --             avalon_slave_L_buffer.address
			avalon_slave_L_buffer_waitrequest  => mm_interconnect_10_comm_pedreiro_v1_01_f_avalon_slave_l_buffer_waitrequest,   --                                  .waitrequest
			avalon_slave_L_buffer_write        => mm_interconnect_10_comm_pedreiro_v1_01_f_avalon_slave_l_buffer_write,         --                                  .write
			avalon_slave_L_buffer_writedata    => mm_interconnect_10_comm_pedreiro_v1_01_f_avalon_slave_l_buffer_writedata,     --                                  .writedata
			avalon_slave_R_buffer_address      => mm_interconnect_16_comm_pedreiro_v1_01_f_avalon_slave_r_buffer_address,       --             avalon_slave_R_buffer.address
			avalon_slave_R_buffer_write        => mm_interconnect_16_comm_pedreiro_v1_01_f_avalon_slave_r_buffer_write,         --                                  .write
			avalon_slave_R_buffer_writedata    => mm_interconnect_16_comm_pedreiro_v1_01_f_avalon_slave_r_buffer_writedata,     --                                  .writedata
			avalon_slave_R_buffer_waitrequest  => mm_interconnect_16_comm_pedreiro_v1_01_f_avalon_slave_r_buffer_waitrequest,   --                                  .waitrequest
			measurements_channel               => comm_f_measurements_conduit_end_measurements_channel_signal,                  --          measurements_conduit_end.measurements_channel_signal
			fee_codec_rmap_wr_waitrequest_i    => rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal,      -- conduit_end_fee_rmap_master_codec.wr_waitrequest_signal
			fee_codec_rmap_readdata_i          => rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_readdata_signal,            --                                  .readdata_signal
			fee_codec_rmap_rd_waitrequest_i    => rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal,      --                                  .rd_waitrequest_signal
			fee_codec_rmap_wr_address_o        => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_wr_address_signal,    --                                  .wr_address_signal
			fee_codec_rmap_write_o             => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_write_signal,         --                                  .write_signal
			fee_codec_rmap_writedata_o         => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_writedata_signal,     --                                  .writedata_signal
			fee_codec_rmap_rd_address_o        => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_rd_address_signal,    --                                  .rd_address_signal
			fee_codec_rmap_read_o              => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_read_signal,          --                                  .read_signal
			fee_hk_rmap_wr_waitrequest_i       => rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal,      --    conduit_end_fee_rmap_master_hk.wr_waitrequest_signal
			fee_hk_rmap_readdata_i             => rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_readdata_signal,            --                                  .readdata_signal
			fee_hk_rmap_rd_waitrequest_i       => rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal,      --                                  .rd_waitrequest_signal
			fee_hk_rmap_wr_address_o           => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_wr_address_signal,       --                                  .wr_address_signal
			fee_hk_rmap_write_o                => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_write_signal,            --                                  .write_signal
			fee_hk_rmap_writedata_o            => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_writedata_signal,        --                                  .writedata_signal
			fee_hk_rmap_rd_address_o           => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_rd_address_signal,       --                                  .rd_address_signal
			fee_hk_rmap_read_o                 => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_read_signal,             --                                  .read_signal
			channel_hk_timecode_control_o      => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_timecode_control_signal,     --        conduit_end_channel_hk_out.timecode_control_signal
			channel_hk_timecode_time_o         => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_timecode_time_signal,        --                                  .timecode_time_signal
			channel_hk_rmap_target_status_o    => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_rmap_target_status_signal,   --                                  .rmap_target_status_signal
			channel_hk_rmap_target_indicate_o  => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_rmap_target_indicate_signal, --                                  .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_o   => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_escape_err_signal,  --                                  .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_o   => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_credit_err_signal,  --                                  .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_o   => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_parity_err_signal,  --                                  .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_o   => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_disconnect_signal,  --                                  .spw_link_disconnect_signal
			channel_hk_spw_link_running_o      => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_running_signal,     --                                  .spw_link_running_signal
			channel_hk_frame_counter_o         => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_frame_counter_signal,        --                                  .frame_counter_signal
			channel_hk_frame_number_o          => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_frame_number_signal,         --                                  .frame_number_signal
			channel_win_mem_addr_offset_o      => comm_pedreiro_v1_01_f_conduit_end_avm_configs_out_win_mem_addr_offset_signal  --       conduit_end_avm_configs_out.win_mem_addr_offset_signal
		);

	ftdi_usb3_0 : component ftdi_usb3_top
		port map (
			clock_sink_clk                  => m2_ddr2_memory_afi_half_clk_clk,                               --            clock_sink.clk
			ftdi_clock_sink_clk             => ftdi_clk_clk,                                                  --       ftdi_clock_sink.clk
			reset_sink_reset                => rst_controller_008_reset_out_reset,                            --            reset_sink.reset
			umft_data_bus                   => umft601a_pins_umft_data_signal,                                --     conduit_umft_pins.umft_data_signal
			umft_reset_n_pin                => umft601a_pins_umft_reset_n_signal,                             --                      .umft_reset_n_signal
			umft_rxf_n_pin                  => umft601a_pins_umft_rxf_n_signal,                               --                      .umft_rxf_n_signal
			umft_clock_pin                  => umft601a_pins_umft_clock_signal,                               --                      .umft_clock_signal
			umft_wakeup_n_pin               => umft601a_pins_umft_wakeup_n_signal,                            --                      .umft_wakeup_n_signal
			umft_be_bus                     => umft601a_pins_umft_be_signal,                                  --                      .umft_be_signal
			umft_txe_n_pin                  => umft601a_pins_umft_txe_n_signal,                               --                      .umft_txe_n_signal
			umft_gpio_bus                   => umft601a_pins_umft_gpio_bus_signal,                            --                      .umft_gpio_bus_signal
			umft_wr_n_pin                   => umft601a_pins_umft_wr_n_signal,                                --                      .umft_wr_n_signal
			umft_rd_n_pin                   => umft601a_pins_umft_rd_n_signal,                                --                      .umft_rd_n_signal
			umft_oe_n_pin                   => umft601a_pins_umft_oe_n_signal,                                --                      .umft_oe_n_signal
			umft_siwu_n_pin                 => umft601a_pins_umft_siwu_n_signal,                              --                      .umft_siwu_n_signal
			avalon_slave_config_address     => mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_address,     --   avalon_slave_config.address
			avalon_slave_config_write       => mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_write,       --                      .write
			avalon_slave_config_read        => mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_read,        --                      .read
			avalon_slave_config_readdata    => mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_readdata,    --                      .readdata
			avalon_slave_config_writedata   => mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_writedata,   --                      .writedata
			avalon_slave_config_waitrequest => mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_waitrequest, --                      .waitrequest
			avalon_slave_config_byteenable  => mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_byteenable,  --                      .byteenable
			avalon_slave_data_address       => mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_address,       --     avalon_slave_data.address
			avalon_slave_data_write         => mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_write,         --                      .write
			avalon_slave_data_read          => mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_read,          --                      .read
			avalon_slave_data_writedata     => mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_writedata,     --                      .writedata
			avalon_slave_data_readdata      => mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_readdata,      --                      .readdata
			avalon_slave_data_waitrequest   => mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_waitrequest,   --                      .waitrequest
			ftdi_interrupt_sender_irq       => irq_mapper_receiver19_irq                                      -- ftdi_interrupt_sender.irq
		);

	seven_segment_controller_0 : component SEVEN_SEG_TOP
		port map (
			AVALON_SLAVE_ADDRESS   => mm_interconnect_2_seven_segment_controller_0_ssdp_avalon_slave_address(0), -- SSDP_avalon_slave.address
			AVALON_SLAVE_WRITEDATA => mm_interconnect_2_seven_segment_controller_0_ssdp_avalon_slave_writedata,  --                  .writedata
			AVALON_SLAVE_WRITE     => mm_interconnect_2_seven_segment_controller_0_ssdp_avalon_slave_write,      --                  .write
			CLK                    => clk50_clk,                                                                 --          SSDP_CLK.clk
			RST                    => rst_controller_009_reset_out_reset,                                        --          SSDP_RST.reset
			SEVEN_SEG_DSP0_OUT     => ssdp_ssdp0,                                                                --      SSDP_conduit.ssdp0
			SEVEN_SEG_DSP1_OUT     => ssdp_ssdp1                                                                 --                  .ssdp1
		);

	clock_bridge_afi_50 : component mebx_qsys_project_clock_bridge_afi_50
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			HDL_ADDR_WIDTH      => 12,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 4,
			RESPONSE_FIFO_DEPTH => 4,
			MASTER_SYNC_DEPTH   => 2,
			SLAVE_SYNC_DEPTH    => 2
		)
		port map (
			m0_clk           => clk50_clk,                                              --   m0_clk.clk
			m0_reset         => rst_controller_009_reset_out_reset,                     -- m0_reset.reset
			s0_clk           => m2_ddr2_memory_afi_half_clk_clk,                        --   s0_clk.clk
			s0_reset         => rst_controller_008_reset_out_reset,                     -- s0_reset.reset
			s0_waitrequest   => mm_interconnect_1_clock_bridge_afi_50_s0_waitrequest,   --       s0.waitrequest
			s0_readdata      => mm_interconnect_1_clock_bridge_afi_50_s0_readdata,      --         .readdata
			s0_readdatavalid => mm_interconnect_1_clock_bridge_afi_50_s0_readdatavalid, --         .readdatavalid
			s0_burstcount    => mm_interconnect_1_clock_bridge_afi_50_s0_burstcount,    --         .burstcount
			s0_writedata     => mm_interconnect_1_clock_bridge_afi_50_s0_writedata,     --         .writedata
			s0_address       => mm_interconnect_1_clock_bridge_afi_50_s0_address,       --         .address
			s0_write         => mm_interconnect_1_clock_bridge_afi_50_s0_write,         --         .write
			s0_read          => mm_interconnect_1_clock_bridge_afi_50_s0_read,          --         .read
			s0_byteenable    => mm_interconnect_1_clock_bridge_afi_50_s0_byteenable,    --         .byteenable
			s0_debugaccess   => mm_interconnect_1_clock_bridge_afi_50_s0_debugaccess,   --         .debugaccess
			m0_waitrequest   => clock_bridge_afi_50_m0_waitrequest,                     --       m0.waitrequest
			m0_readdata      => clock_bridge_afi_50_m0_readdata,                        --         .readdata
			m0_readdatavalid => clock_bridge_afi_50_m0_readdatavalid,                   --         .readdatavalid
			m0_burstcount    => clock_bridge_afi_50_m0_burstcount,                      --         .burstcount
			m0_writedata     => clock_bridge_afi_50_m0_writedata,                       --         .writedata
			m0_address       => clock_bridge_afi_50_m0_address,                         --         .address
			m0_write         => clock_bridge_afi_50_m0_write,                           --         .write
			m0_read          => clock_bridge_afi_50_m0_read,                            --         .read
			m0_byteenable    => clock_bridge_afi_50_m0_byteenable,                      --         .byteenable
			m0_debugaccess   => clock_bridge_afi_50_m0_debugaccess                      --         .debugaccess
		);

	csense_adc_fo : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                          --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_2_csense_adc_fo_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_csense_adc_fo_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_csense_adc_fo_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_csense_adc_fo_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_csense_adc_fo_s1_readdata,        --                    .readdata
			out_port   => csense_adc_fo_export                                -- external_connection.export
		);

	csense_cs_n : component MebX_Qsys_Project_csense_cs_n
		port map (
			clk        => clk50_clk,                                        --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_2_csense_cs_n_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_csense_cs_n_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_csense_cs_n_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_csense_cs_n_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_csense_cs_n_s1_readdata,        --                    .readdata
			out_port   => csense_cs_n_export                                -- external_connection.export
		);

	csense_sck : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                       --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_2_csense_sck_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_csense_sck_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_csense_sck_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_csense_sck_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_csense_sck_s1_readdata,        --                    .readdata
			out_port   => csense_sck_export                                -- external_connection.export
		);

	csense_sdi : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                       --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_2_csense_sdi_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_csense_sdi_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_csense_sdi_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_csense_sdi_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_csense_sdi_s1_readdata,        --                    .readdata
			out_port   => csense_sdi_export                                -- external_connection.export
		);

	csense_sdo : component MebX_Qsys_Project_csense_sdo
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_009_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_csense_sdo_s1_address,      --                  s1.address
			readdata => mm_interconnect_2_csense_sdo_s1_readdata,     --                    .readdata
			in_port  => csense_sdo_export                             -- external_connection.export
		);

	ddr2_address_span_extender : component altera_address_span_extender
		generic map (
			DATA_WIDTH           => 32,
			BYTEENABLE_WIDTH     => 4,
			MASTER_ADDRESS_WIDTH => 32,
			SLAVE_ADDRESS_WIDTH  => 29,
			SLAVE_ADDRESS_SHIFT  => 2,
			BURSTCOUNT_WIDTH     => 8,
			CNTL_ADDRESS_WIDTH   => 1,
			SUB_WINDOW_COUNT     => 1,
			MASTER_ADDRESS_DEF   => "0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			clk                  => m2_ddr2_memory_afi_half_clk_clk,                                           --           clock.clk
			reset                => rst_controller_008_reset_out_reset,                                        --           reset.reset
			avs_s0_address       => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_address,       --  windowed_slave.address
			avs_s0_read          => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_read,          --                .read
			avs_s0_readdata      => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdata,      --                .readdata
			avs_s0_write         => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_write,         --                .write
			avs_s0_writedata     => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_writedata,     --                .writedata
			avs_s0_readdatavalid => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdatavalid, --                .readdatavalid
			avs_s0_waitrequest   => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_waitrequest,   --                .waitrequest
			avs_s0_byteenable    => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_byteenable,    --                .byteenable
			avs_s0_burstcount    => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_burstcount,    --                .burstcount
			avm_m0_address       => ddr2_address_span_extender_expanded_master_address,                        -- expanded_master.address
			avm_m0_read          => ddr2_address_span_extender_expanded_master_read,                           --                .read
			avm_m0_waitrequest   => ddr2_address_span_extender_expanded_master_waitrequest,                    --                .waitrequest
			avm_m0_readdata      => ddr2_address_span_extender_expanded_master_readdata,                       --                .readdata
			avm_m0_write         => ddr2_address_span_extender_expanded_master_write,                          --                .write
			avm_m0_writedata     => ddr2_address_span_extender_expanded_master_writedata,                      --                .writedata
			avm_m0_readdatavalid => ddr2_address_span_extender_expanded_master_readdatavalid,                  --                .readdatavalid
			avm_m0_byteenable    => ddr2_address_span_extender_expanded_master_byteenable,                     --                .byteenable
			avm_m0_burstcount    => ddr2_address_span_extender_expanded_master_burstcount,                     --                .burstcount
			avs_cntl_read        => mm_interconnect_1_ddr2_address_span_extender_cntl_read,                    --            cntl.read
			avs_cntl_readdata    => mm_interconnect_1_ddr2_address_span_extender_cntl_readdata,                --                .readdata
			avs_cntl_write       => mm_interconnect_1_ddr2_address_span_extender_cntl_write,                   --                .write
			avs_cntl_writedata   => mm_interconnect_1_ddr2_address_span_extender_cntl_writedata,               --                .writedata
			avs_cntl_byteenable  => mm_interconnect_1_ddr2_address_span_extender_cntl_byteenable,              --                .byteenable
			avs_cntl_address     => "0"                                                                        --     (terminated)
		);

	dma_comm_1_left : component MebX_Qsys_Project_dma_comm_1_left
		port map (
			mm_read_address              => dma_comm_1_left_mm_read_address,                                --          mm_read.address
			mm_read_read                 => dma_comm_1_left_mm_read_read,                                   --                 .read
			mm_read_byteenable           => dma_comm_1_left_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => dma_comm_1_left_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => dma_comm_1_left_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => dma_comm_1_left_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_write_address             => dma_comm_1_left_mm_write_address,                               --         mm_write.address
			mm_write_write               => dma_comm_1_left_mm_write_write,                                 --                 .write
			mm_write_byteenable          => dma_comm_1_left_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => dma_comm_1_left_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => dma_comm_1_left_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => m2_ddr2_memory_afi_half_clk_clk,                                --            clock.clk
			reset_n_reset_n              => rst_controller_008_reset_out_reset_ports_inv,                   --          reset_n.reset_n
			csr_writedata                => mm_interconnect_1_dma_comm_1_left_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_1_dma_comm_1_left_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_1_dma_comm_1_left_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_1_dma_comm_1_left_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_1_dma_comm_1_left_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_1_dma_comm_1_left_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_1_dma_comm_1_left_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_1_dma_comm_1_left_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_1_dma_comm_1_left_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_1_dma_comm_1_left_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver6_irq                                        --          csr_irq.irq
		);

	dma_comm_1_right : component MebX_Qsys_Project_dma_comm_1_right
		port map (
			mm_read_address              => dma_comm_1_right_mm_read_address,                                --          mm_read.address
			mm_read_read                 => dma_comm_1_right_mm_read_read,                                   --                 .read
			mm_read_byteenable           => dma_comm_1_right_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => dma_comm_1_right_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => dma_comm_1_right_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => dma_comm_1_right_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_write_address             => dma_comm_1_right_mm_write_address,                               --         mm_write.address
			mm_write_write               => dma_comm_1_right_mm_write_write,                                 --                 .write
			mm_write_byteenable          => dma_comm_1_right_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => dma_comm_1_right_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => dma_comm_1_right_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => m2_ddr2_memory_afi_half_clk_clk,                                 --            clock.clk
			reset_n_reset_n              => rst_controller_008_reset_out_reset_ports_inv,                    --          reset_n.reset_n
			csr_writedata                => mm_interconnect_1_dma_comm_1_right_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_1_dma_comm_1_right_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_1_dma_comm_1_right_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_1_dma_comm_1_right_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_1_dma_comm_1_right_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_1_dma_comm_1_right_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_1_dma_comm_1_right_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_1_dma_comm_1_right_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_1_dma_comm_1_right_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_1_dma_comm_1_right_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver7_irq                                         --          csr_irq.irq
		);

	dma_comm_2_left : component MebX_Qsys_Project_dma_comm_2_left
		port map (
			mm_read_address              => dma_comm_2_left_mm_read_address,                                --          mm_read.address
			mm_read_read                 => dma_comm_2_left_mm_read_read,                                   --                 .read
			mm_read_byteenable           => dma_comm_2_left_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => dma_comm_2_left_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => dma_comm_2_left_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => dma_comm_2_left_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_write_address             => dma_comm_2_left_mm_write_address,                               --         mm_write.address
			mm_write_write               => dma_comm_2_left_mm_write_write,                                 --                 .write
			mm_write_byteenable          => dma_comm_2_left_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => dma_comm_2_left_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => dma_comm_2_left_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => m2_ddr2_memory_afi_half_clk_clk,                                --            clock.clk
			reset_n_reset_n              => rst_controller_008_reset_out_reset_ports_inv,                   --          reset_n.reset_n
			csr_writedata                => mm_interconnect_1_dma_comm_2_left_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_1_dma_comm_2_left_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_1_dma_comm_2_left_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_1_dma_comm_2_left_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_1_dma_comm_2_left_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_1_dma_comm_2_left_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_1_dma_comm_2_left_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_1_dma_comm_2_left_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_1_dma_comm_2_left_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_1_dma_comm_2_left_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver8_irq                                        --          csr_irq.irq
		);

	dma_comm_2_right : component MebX_Qsys_Project_dma_comm_2_right
		port map (
			mm_read_address              => dma_comm_2_right_mm_read_address,                                --          mm_read.address
			mm_read_read                 => dma_comm_2_right_mm_read_read,                                   --                 .read
			mm_read_byteenable           => dma_comm_2_right_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => dma_comm_2_right_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => dma_comm_2_right_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => dma_comm_2_right_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_write_address             => dma_comm_2_right_mm_write_address,                               --         mm_write.address
			mm_write_write               => dma_comm_2_right_mm_write_write,                                 --                 .write
			mm_write_byteenable          => dma_comm_2_right_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => dma_comm_2_right_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => dma_comm_2_right_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => m2_ddr2_memory_afi_half_clk_clk,                                 --            clock.clk
			reset_n_reset_n              => rst_controller_008_reset_out_reset_ports_inv,                    --          reset_n.reset_n
			csr_writedata                => mm_interconnect_1_dma_comm_2_right_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_1_dma_comm_2_right_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_1_dma_comm_2_right_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_1_dma_comm_2_right_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_1_dma_comm_2_right_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_1_dma_comm_2_right_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_1_dma_comm_2_right_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_1_dma_comm_2_right_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_1_dma_comm_2_right_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_1_dma_comm_2_right_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver9_irq                                         --          csr_irq.irq
		);

	dma_comm_3_left : component MebX_Qsys_Project_dma_comm_3_left
		port map (
			mm_read_address              => dma_comm_3_left_mm_read_address,                                --          mm_read.address
			mm_read_read                 => dma_comm_3_left_mm_read_read,                                   --                 .read
			mm_read_byteenable           => dma_comm_3_left_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => dma_comm_3_left_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => dma_comm_3_left_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => dma_comm_3_left_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_write_address             => dma_comm_3_left_mm_write_address,                               --         mm_write.address
			mm_write_write               => dma_comm_3_left_mm_write_write,                                 --                 .write
			mm_write_byteenable          => dma_comm_3_left_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => dma_comm_3_left_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => dma_comm_3_left_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => m2_ddr2_memory_afi_half_clk_clk,                                --            clock.clk
			reset_n_reset_n              => rst_controller_008_reset_out_reset_ports_inv,                   --          reset_n.reset_n
			csr_writedata                => mm_interconnect_1_dma_comm_3_left_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_1_dma_comm_3_left_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_1_dma_comm_3_left_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_1_dma_comm_3_left_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_1_dma_comm_3_left_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_1_dma_comm_3_left_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_1_dma_comm_3_left_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_1_dma_comm_3_left_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_1_dma_comm_3_left_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_1_dma_comm_3_left_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver10_irq                                       --          csr_irq.irq
		);

	dma_comm_3_right : component MebX_Qsys_Project_dma_comm_3_right
		port map (
			mm_read_address              => dma_comm_3_right_mm_read_address,                                --          mm_read.address
			mm_read_read                 => dma_comm_3_right_mm_read_read,                                   --                 .read
			mm_read_byteenable           => dma_comm_3_right_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => dma_comm_3_right_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => dma_comm_3_right_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => dma_comm_3_right_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_write_address             => dma_comm_3_right_mm_write_address,                               --         mm_write.address
			mm_write_write               => dma_comm_3_right_mm_write_write,                                 --                 .write
			mm_write_byteenable          => dma_comm_3_right_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => dma_comm_3_right_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => dma_comm_3_right_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => m2_ddr2_memory_afi_half_clk_clk,                                 --            clock.clk
			reset_n_reset_n              => rst_controller_008_reset_out_reset_ports_inv,                    --          reset_n.reset_n
			csr_writedata                => mm_interconnect_1_dma_comm_3_right_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_1_dma_comm_3_right_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_1_dma_comm_3_right_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_1_dma_comm_3_right_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_1_dma_comm_3_right_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_1_dma_comm_3_right_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_1_dma_comm_3_right_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_1_dma_comm_3_right_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_1_dma_comm_3_right_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_1_dma_comm_3_right_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver11_irq                                        --          csr_irq.irq
		);

	dma_comm_4_left : component MebX_Qsys_Project_dma_comm_4_left
		port map (
			mm_read_address              => dma_comm_4_left_mm_read_address,                                --          mm_read.address
			mm_read_read                 => dma_comm_4_left_mm_read_read,                                   --                 .read
			mm_read_byteenable           => dma_comm_4_left_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => dma_comm_4_left_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => dma_comm_4_left_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => dma_comm_4_left_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_write_address             => dma_comm_4_left_mm_write_address,                               --         mm_write.address
			mm_write_write               => dma_comm_4_left_mm_write_write,                                 --                 .write
			mm_write_byteenable          => dma_comm_4_left_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => dma_comm_4_left_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => dma_comm_4_left_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => m2_ddr2_memory_afi_half_clk_clk,                                --            clock.clk
			reset_n_reset_n              => rst_controller_008_reset_out_reset_ports_inv,                   --          reset_n.reset_n
			csr_writedata                => mm_interconnect_1_dma_comm_4_left_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_1_dma_comm_4_left_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_1_dma_comm_4_left_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_1_dma_comm_4_left_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_1_dma_comm_4_left_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_1_dma_comm_4_left_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_1_dma_comm_4_left_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_1_dma_comm_4_left_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_1_dma_comm_4_left_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_1_dma_comm_4_left_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver12_irq                                       --          csr_irq.irq
		);

	dma_comm_4_right : component MebX_Qsys_Project_dma_comm_4_right
		port map (
			mm_read_address              => dma_comm_4_right_mm_read_address,                                --          mm_read.address
			mm_read_read                 => dma_comm_4_right_mm_read_read,                                   --                 .read
			mm_read_byteenable           => dma_comm_4_right_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => dma_comm_4_right_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => dma_comm_4_right_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => dma_comm_4_right_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_write_address             => dma_comm_4_right_mm_write_address,                               --         mm_write.address
			mm_write_write               => dma_comm_4_right_mm_write_write,                                 --                 .write
			mm_write_byteenable          => dma_comm_4_right_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => dma_comm_4_right_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => dma_comm_4_right_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => m2_ddr2_memory_afi_half_clk_clk,                                 --            clock.clk
			reset_n_reset_n              => rst_controller_008_reset_out_reset_ports_inv,                    --          reset_n.reset_n
			csr_writedata                => mm_interconnect_1_dma_comm_4_right_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_1_dma_comm_4_right_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_1_dma_comm_4_right_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_1_dma_comm_4_right_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_1_dma_comm_4_right_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_1_dma_comm_4_right_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_1_dma_comm_4_right_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_1_dma_comm_4_right_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_1_dma_comm_4_right_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_1_dma_comm_4_right_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver13_irq                                        --          csr_irq.irq
		);

	dma_comm_5_left : component MebX_Qsys_Project_dma_comm_5_left
		port map (
			mm_read_address              => dma_comm_5_left_mm_read_address,                                --          mm_read.address
			mm_read_read                 => dma_comm_5_left_mm_read_read,                                   --                 .read
			mm_read_byteenable           => dma_comm_5_left_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => dma_comm_5_left_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => dma_comm_5_left_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => dma_comm_5_left_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_write_address             => dma_comm_5_left_mm_write_address,                               --         mm_write.address
			mm_write_write               => dma_comm_5_left_mm_write_write,                                 --                 .write
			mm_write_byteenable          => dma_comm_5_left_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => dma_comm_5_left_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => dma_comm_5_left_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => m2_ddr2_memory_afi_half_clk_clk,                                --            clock.clk
			reset_n_reset_n              => rst_controller_008_reset_out_reset_ports_inv,                   --          reset_n.reset_n
			csr_writedata                => mm_interconnect_1_dma_comm_5_left_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_1_dma_comm_5_left_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_1_dma_comm_5_left_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_1_dma_comm_5_left_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_1_dma_comm_5_left_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_1_dma_comm_5_left_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_1_dma_comm_5_left_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_1_dma_comm_5_left_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_1_dma_comm_5_left_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_1_dma_comm_5_left_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver17_irq                                       --          csr_irq.irq
		);

	dma_comm_5_right : component MebX_Qsys_Project_dma_comm_5_right
		port map (
			mm_read_address              => dma_comm_5_right_mm_read_address,                                --          mm_read.address
			mm_read_read                 => dma_comm_5_right_mm_read_read,                                   --                 .read
			mm_read_byteenable           => dma_comm_5_right_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => dma_comm_5_right_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => dma_comm_5_right_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => dma_comm_5_right_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_write_address             => dma_comm_5_right_mm_write_address,                               --         mm_write.address
			mm_write_write               => dma_comm_5_right_mm_write_write,                                 --                 .write
			mm_write_byteenable          => dma_comm_5_right_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => dma_comm_5_right_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => dma_comm_5_right_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => m2_ddr2_memory_afi_half_clk_clk,                                 --            clock.clk
			reset_n_reset_n              => rst_controller_008_reset_out_reset_ports_inv,                    --          reset_n.reset_n
			csr_writedata                => mm_interconnect_1_dma_comm_5_right_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_1_dma_comm_5_right_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_1_dma_comm_5_right_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_1_dma_comm_5_right_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_1_dma_comm_5_right_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_1_dma_comm_5_right_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_1_dma_comm_5_right_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_1_dma_comm_5_right_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_1_dma_comm_5_right_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_1_dma_comm_5_right_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver16_irq                                        --          csr_irq.irq
		);

	dma_comm_6_left : component MebX_Qsys_Project_dma_comm_6_left
		port map (
			mm_read_address              => dma_comm_6_left_mm_read_address,                                --          mm_read.address
			mm_read_read                 => dma_comm_6_left_mm_read_read,                                   --                 .read
			mm_read_byteenable           => dma_comm_6_left_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => dma_comm_6_left_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => dma_comm_6_left_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => dma_comm_6_left_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_write_address             => dma_comm_6_left_mm_write_address,                               --         mm_write.address
			mm_write_write               => dma_comm_6_left_mm_write_write,                                 --                 .write
			mm_write_byteenable          => dma_comm_6_left_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => dma_comm_6_left_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => dma_comm_6_left_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => m2_ddr2_memory_afi_half_clk_clk,                                --            clock.clk
			reset_n_reset_n              => rst_controller_008_reset_out_reset_ports_inv,                   --          reset_n.reset_n
			csr_writedata                => mm_interconnect_1_dma_comm_6_left_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_1_dma_comm_6_left_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_1_dma_comm_6_left_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_1_dma_comm_6_left_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_1_dma_comm_6_left_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_1_dma_comm_6_left_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_1_dma_comm_6_left_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_1_dma_comm_6_left_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_1_dma_comm_6_left_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_1_dma_comm_6_left_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver15_irq                                       --          csr_irq.irq
		);

	dma_comm_6_right : component MebX_Qsys_Project_dma_comm_6_right
		port map (
			mm_read_address              => dma_comm_6_right_mm_read_address,                                --          mm_read.address
			mm_read_read                 => dma_comm_6_right_mm_read_read,                                   --                 .read
			mm_read_byteenable           => dma_comm_6_right_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => dma_comm_6_right_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => dma_comm_6_right_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => dma_comm_6_right_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_write_address             => dma_comm_6_right_mm_write_address,                               --         mm_write.address
			mm_write_write               => dma_comm_6_right_mm_write_write,                                 --                 .write
			mm_write_byteenable          => dma_comm_6_right_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => dma_comm_6_right_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => dma_comm_6_right_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => m2_ddr2_memory_afi_half_clk_clk,                                 --            clock.clk
			reset_n_reset_n              => rst_controller_008_reset_out_reset_ports_inv,                    --          reset_n.reset_n
			csr_writedata                => mm_interconnect_1_dma_comm_6_right_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_1_dma_comm_6_right_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_1_dma_comm_6_right_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_1_dma_comm_6_right_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_1_dma_comm_6_right_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_1_dma_comm_6_right_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_1_dma_comm_6_right_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_1_dma_comm_6_right_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_1_dma_comm_6_right_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_1_dma_comm_6_right_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver14_irq                                        --          csr_irq.irq
		);

	dma_ftdi_usb3 : component MebX_Qsys_Project_dma_ftdi_usb3
		port map (
			mm_read_address              => dma_ftdi_usb3_mm_read_address,                                --          mm_read.address
			mm_read_read                 => dma_ftdi_usb3_mm_read_read,                                   --                 .read
			mm_read_byteenable           => dma_ftdi_usb3_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => dma_ftdi_usb3_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => dma_ftdi_usb3_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => dma_ftdi_usb3_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_write_address             => dma_ftdi_usb3_mm_write_address,                               --         mm_write.address
			mm_write_write               => dma_ftdi_usb3_mm_write_write,                                 --                 .write
			mm_write_byteenable          => dma_ftdi_usb3_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => dma_ftdi_usb3_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => dma_ftdi_usb3_mm_write_waitrequest,                           --                 .waitrequest
			clock_clk                    => m2_ddr2_memory_afi_half_clk_clk,                              --            clock.clk
			reset_n_reset_n              => rst_controller_008_reset_out_reset_ports_inv,                 --          reset_n.reset_n
			csr_writedata                => mm_interconnect_1_dma_ftdi_usb3_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_1_dma_ftdi_usb3_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_1_dma_ftdi_usb3_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_1_dma_ftdi_usb3_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_1_dma_ftdi_usb3_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_1_dma_ftdi_usb3_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_1_dma_ftdi_usb3_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_1_dma_ftdi_usb3_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_1_dma_ftdi_usb3_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_1_dma_ftdi_usb3_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver18_irq                                     --          csr_irq.irq
		);

	ext_flash : component MebX_Qsys_Project_ext_flash
		generic map (
			TCM_ADDRESS_W                  => 26,
			TCM_DATA_W                     => 16,
			TCM_BYTEENABLE_W               => 2,
			TCM_READ_WAIT                  => 100,
			TCM_WRITE_WAIT                 => 100,
			TCM_SETUP_WAIT                 => 25,
			TCM_DATA_HOLD                  => 20,
			TCM_TURNAROUND_TIME            => 2,
			TCM_TIMING_UNITS               => 0,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 2,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 1,
			USE_WRITE                      => 1,
			USE_BYTEENABLE                 => 0,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 0,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 0,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 0,
			ACTIVE_LOW_READ                => 1,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 1,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 0,
			ACTIVE_LOW_OUTPUTENABLE        => 0,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0
		)
		port map (
			clk_clk              => m2_ddr2_memory_afi_half_clk_clk,               --   clk.clk
			reset_reset          => rst_controller_010_reset_out_reset,            -- reset.reset
			uas_address          => mm_interconnect_1_ext_flash_uas_address,       --   uas.address
			uas_burstcount       => mm_interconnect_1_ext_flash_uas_burstcount,    --      .burstcount
			uas_read             => mm_interconnect_1_ext_flash_uas_read,          --      .read
			uas_write            => mm_interconnect_1_ext_flash_uas_write,         --      .write
			uas_waitrequest      => mm_interconnect_1_ext_flash_uas_waitrequest,   --      .waitrequest
			uas_readdatavalid    => mm_interconnect_1_ext_flash_uas_readdatavalid, --      .readdatavalid
			uas_byteenable       => mm_interconnect_1_ext_flash_uas_byteenable,    --      .byteenable
			uas_readdata         => mm_interconnect_1_ext_flash_uas_readdata,      --      .readdata
			uas_writedata        => mm_interconnect_1_ext_flash_uas_writedata,     --      .writedata
			uas_lock             => mm_interconnect_1_ext_flash_uas_lock,          --      .lock
			uas_debugaccess      => mm_interconnect_1_ext_flash_uas_debugaccess,   --      .debugaccess
			tcm_write_n_out      => ext_flash_tcm_write_n_out,                     --   tcm.write_n_out
			tcm_read_n_out       => ext_flash_tcm_read_n_out,                      --      .read_n_out
			tcm_chipselect_n_out => ext_flash_tcm_chipselect_n_out,                --      .chipselect_n_out
			tcm_request          => ext_flash_tcm_request,                         --      .request
			tcm_grant            => ext_flash_tcm_grant,                           --      .grant
			tcm_address_out      => ext_flash_tcm_address_out,                     --      .address_out
			tcm_data_out         => ext_flash_tcm_data_out,                        --      .data_out
			tcm_data_outen       => ext_flash_tcm_data_outen,                      --      .data_outen
			tcm_data_in          => ext_flash_tcm_data_in                          --      .data_in
		);

	jtag_uart_0 : component MebX_Qsys_Project_jtag_uart_0
		port map (
			clk            => m2_ddr2_memory_afi_half_clk_clk,                                 --               clk.clk
			rst_n          => rst_controller_008_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver20_irq                                        --               irq.irq
		);

	m1_clock_bridge : component mebx_qsys_project_m1_clock_bridge
		generic map (
			DATA_WIDTH          => 256,
			SYMBOL_WIDTH        => 8,
			HDL_ADDR_WIDTH      => 31,
			BURSTCOUNT_WIDTH    => 3,
			COMMAND_FIFO_DEPTH  => 8,
			RESPONSE_FIFO_DEPTH => 8,
			MASTER_SYNC_DEPTH   => 2,
			SLAVE_SYNC_DEPTH    => 2
		)
		port map (
			m0_clk           => m1_ddr2_memory_afi_half_clk_clk,                    --   m0_clk.clk
			m0_reset         => rst_controller_011_reset_out_reset,                 -- m0_reset.reset
			s0_clk           => m2_ddr2_memory_afi_half_clk_clk,                    --   s0_clk.clk
			s0_reset         => rst_controller_008_reset_out_reset,                 -- s0_reset.reset
			s0_waitrequest   => mm_interconnect_0_m1_clock_bridge_s0_waitrequest,   --       s0.waitrequest
			s0_readdata      => mm_interconnect_0_m1_clock_bridge_s0_readdata,      --         .readdata
			s0_readdatavalid => mm_interconnect_0_m1_clock_bridge_s0_readdatavalid, --         .readdatavalid
			s0_burstcount    => mm_interconnect_0_m1_clock_bridge_s0_burstcount,    --         .burstcount
			s0_writedata     => mm_interconnect_0_m1_clock_bridge_s0_writedata,     --         .writedata
			s0_address       => mm_interconnect_0_m1_clock_bridge_s0_address,       --         .address
			s0_write         => mm_interconnect_0_m1_clock_bridge_s0_write,         --         .write
			s0_read          => mm_interconnect_0_m1_clock_bridge_s0_read,          --         .read
			s0_byteenable    => mm_interconnect_0_m1_clock_bridge_s0_byteenable,    --         .byteenable
			s0_debugaccess   => mm_interconnect_0_m1_clock_bridge_s0_debugaccess,   --         .debugaccess
			m0_waitrequest   => m1_clock_bridge_m0_waitrequest,                     --       m0.waitrequest
			m0_readdata      => m1_clock_bridge_m0_readdata,                        --         .readdata
			m0_readdatavalid => m1_clock_bridge_m0_readdatavalid,                   --         .readdatavalid
			m0_burstcount    => m1_clock_bridge_m0_burstcount,                      --         .burstcount
			m0_writedata     => m1_clock_bridge_m0_writedata,                       --         .writedata
			m0_address       => m1_clock_bridge_m0_address,                         --         .address
			m0_write         => m1_clock_bridge_m0_write,                           --         .write
			m0_read          => m1_clock_bridge_m0_read,                            --         .read
			m0_byteenable    => m1_clock_bridge_m0_byteenable,                      --         .byteenable
			m0_debugaccess   => m1_clock_bridge_m0_debugaccess                      --         .debugaccess
		);

	m1_ddr2_i2c_scl : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                            --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_2_m1_ddr2_i2c_scl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_m1_ddr2_i2c_scl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_m1_ddr2_i2c_scl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_m1_ddr2_i2c_scl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_m1_ddr2_i2c_scl_s1_readdata,        --                    .readdata
			out_port   => m1_ddr2_i2c_scl_export                                -- external_connection.export
		);

	m1_ddr2_i2c_sda : component MebX_Qsys_Project_m1_ddr2_i2c_sda
		port map (
			clk        => clk50_clk,                                            --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_2_m1_ddr2_i2c_sda_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_m1_ddr2_i2c_sda_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_m1_ddr2_i2c_sda_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_m1_ddr2_i2c_sda_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_m1_ddr2_i2c_sda_s1_readdata,        --                    .readdata
			bidir_port => m1_ddr2_i2c_sda_export                                -- external_connection.export
		);

	m1_ddr2_memory : component MebX_Qsys_Project_m1_ddr2_memory
		port map (
			pll_ref_clk        => m1_ddr2_memory_pll_ref_clk_clk,                          --      pll_ref_clk.clk
			global_reset_n     => rst_reset_n,                                             --     global_reset.reset_n
			soft_reset_n       => rst_reset_n,                                             --       soft_reset.reset_n
			afi_clk            => m1_ddr2_memory_afi_clk_clk,                              --          afi_clk.clk
			afi_half_clk       => m1_ddr2_memory_afi_half_clk_clk,                         --     afi_half_clk.clk
			afi_reset_n        => open,                                                    --        afi_reset.reset_n
			afi_reset_export_n => open,                                                    -- afi_reset_export.reset_n
			mem_a              => m1_ddr2_memory_mem_a,                                    --           memory.mem_a
			mem_ba             => m1_ddr2_memory_mem_ba,                                   --                 .mem_ba
			mem_ck             => m1_ddr2_memory_mem_ck,                                   --                 .mem_ck
			mem_ck_n           => m1_ddr2_memory_mem_ck_n,                                 --                 .mem_ck_n
			mem_cke            => m1_ddr2_memory_mem_cke,                                  --                 .mem_cke
			mem_cs_n           => m1_ddr2_memory_mem_cs_n,                                 --                 .mem_cs_n
			mem_dm             => m1_ddr2_memory_mem_dm,                                   --                 .mem_dm
			mem_ras_n          => m1_ddr2_memory_mem_ras_n,                                --                 .mem_ras_n
			mem_cas_n          => m1_ddr2_memory_mem_cas_n,                                --                 .mem_cas_n
			mem_we_n           => m1_ddr2_memory_mem_we_n,                                 --                 .mem_we_n
			mem_dq             => m1_ddr2_memory_mem_dq,                                   --                 .mem_dq
			mem_dqs            => m1_ddr2_memory_mem_dqs,                                  --                 .mem_dqs
			mem_dqs_n          => m1_ddr2_memory_mem_dqs_n,                                --                 .mem_dqs_n
			mem_odt            => m1_ddr2_memory_mem_odt,                                  --                 .mem_odt
			avl_ready          => m1_ddr2_memory_avl_waitrequest,                          --              avl.waitrequest_n
			avl_burstbegin     => mm_interconnect_3_m1_ddr2_memory_avl_beginbursttransfer, --                 .beginbursttransfer
			avl_addr           => mm_interconnect_3_m1_ddr2_memory_avl_address,            --                 .address
			avl_rdata_valid    => mm_interconnect_3_m1_ddr2_memory_avl_readdatavalid,      --                 .readdatavalid
			avl_rdata          => mm_interconnect_3_m1_ddr2_memory_avl_readdata,           --                 .readdata
			avl_wdata          => mm_interconnect_3_m1_ddr2_memory_avl_writedata,          --                 .writedata
			avl_be             => mm_interconnect_3_m1_ddr2_memory_avl_byteenable,         --                 .byteenable
			avl_read_req       => mm_interconnect_3_m1_ddr2_memory_avl_read,               --                 .read
			avl_write_req      => mm_interconnect_3_m1_ddr2_memory_avl_write,              --                 .write
			avl_size           => mm_interconnect_3_m1_ddr2_memory_avl_burstcount,         --                 .burstcount
			local_init_done    => m1_ddr2_memory_status_local_init_done,                   --           status.local_init_done
			local_cal_success  => m1_ddr2_memory_status_local_cal_success,                 --                 .local_cal_success
			local_cal_fail     => m1_ddr2_memory_status_local_cal_fail,                    --                 .local_cal_fail
			oct_rdn            => m1_ddr2_oct_rdn,                                         --              oct.rdn
			oct_rup            => m1_ddr2_oct_rup                                          --                 .rup
		);

	m2_ddr2_i2c_scl : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                            --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_2_m2_ddr2_i2c_scl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_m2_ddr2_i2c_scl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_m2_ddr2_i2c_scl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_m2_ddr2_i2c_scl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_m2_ddr2_i2c_scl_s1_readdata,        --                    .readdata
			out_port   => m2_ddr2_i2c_scl_export                                -- external_connection.export
		);

	m2_ddr2_i2c_sda : component MebX_Qsys_Project_m1_ddr2_i2c_sda
		port map (
			clk        => clk50_clk,                                            --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_2_m2_ddr2_i2c_sda_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_m2_ddr2_i2c_sda_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_m2_ddr2_i2c_sda_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_m2_ddr2_i2c_sda_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_m2_ddr2_i2c_sda_s1_readdata,        --                    .readdata
			bidir_port => m2_ddr2_i2c_sda_export                                -- external_connection.export
		);

	m2_ddr2_memory : component MebX_Qsys_Project_m2_ddr2_memory
		port map (
			pll_ref_clk               => clk50_clk,                                               --      pll_ref_clk.clk
			global_reset_n            => rst_reset_n,                                             --     global_reset.reset_n
			soft_reset_n              => rst_reset_n,                                             --       soft_reset.reset_n
			afi_clk                   => m2_ddr2_memory_afi_clk_clk,                              --          afi_clk.clk
			afi_half_clk              => m2_ddr2_memory_afi_half_clk_clk,                         --     afi_half_clk.clk
			afi_reset_n               => open,                                                    --        afi_reset.reset_n
			afi_reset_export_n        => open,                                                    -- afi_reset_export.reset_n
			mem_a                     => m2_ddr2_memory_mem_a,                                    --           memory.mem_a
			mem_ba                    => m2_ddr2_memory_mem_ba,                                   --                 .mem_ba
			mem_ck                    => m2_ddr2_memory_mem_ck,                                   --                 .mem_ck
			mem_ck_n                  => m2_ddr2_memory_mem_ck_n,                                 --                 .mem_ck_n
			mem_cke                   => m2_ddr2_memory_mem_cke,                                  --                 .mem_cke
			mem_cs_n                  => m2_ddr2_memory_mem_cs_n,                                 --                 .mem_cs_n
			mem_dm                    => m2_ddr2_memory_mem_dm,                                   --                 .mem_dm
			mem_ras_n                 => m2_ddr2_memory_mem_ras_n,                                --                 .mem_ras_n
			mem_cas_n                 => m2_ddr2_memory_mem_cas_n,                                --                 .mem_cas_n
			mem_we_n                  => m2_ddr2_memory_mem_we_n,                                 --                 .mem_we_n
			mem_dq                    => m2_ddr2_memory_mem_dq,                                   --                 .mem_dq
			mem_dqs                   => m2_ddr2_memory_mem_dqs,                                  --                 .mem_dqs
			mem_dqs_n                 => m2_ddr2_memory_mem_dqs_n,                                --                 .mem_dqs_n
			mem_odt                   => m2_ddr2_memory_mem_odt,                                  --                 .mem_odt
			avl_ready                 => m2_ddr2_memory_avl_waitrequest,                          --              avl.waitrequest_n
			avl_burstbegin            => mm_interconnect_0_m2_ddr2_memory_avl_beginbursttransfer, --                 .beginbursttransfer
			avl_addr                  => mm_interconnect_0_m2_ddr2_memory_avl_address,            --                 .address
			avl_rdata_valid           => mm_interconnect_0_m2_ddr2_memory_avl_readdatavalid,      --                 .readdatavalid
			avl_rdata                 => mm_interconnect_0_m2_ddr2_memory_avl_readdata,           --                 .readdata
			avl_wdata                 => mm_interconnect_0_m2_ddr2_memory_avl_writedata,          --                 .writedata
			avl_be                    => mm_interconnect_0_m2_ddr2_memory_avl_byteenable,         --                 .byteenable
			avl_read_req              => mm_interconnect_0_m2_ddr2_memory_avl_read,               --                 .read
			avl_write_req             => mm_interconnect_0_m2_ddr2_memory_avl_write,              --                 .write
			avl_size                  => mm_interconnect_0_m2_ddr2_memory_avl_burstcount,         --                 .burstcount
			local_init_done           => m2_ddr2_memory_status_local_init_done,                   --           status.local_init_done
			local_cal_success         => m2_ddr2_memory_status_local_cal_success,                 --                 .local_cal_success
			local_cal_fail            => m2_ddr2_memory_status_local_cal_fail,                    --                 .local_cal_fail
			oct_rdn                   => m2_ddr2_oct_rdn,                                         --              oct.rdn
			oct_rup                   => m2_ddr2_oct_rup,                                         --                 .rup
			pll_mem_clk               => m2_ddr2_memory_pll_sharing_pll_mem_clk,                  --      pll_sharing.pll_mem_clk
			pll_write_clk             => m2_ddr2_memory_pll_sharing_pll_write_clk,                --                 .pll_write_clk
			pll_locked                => m2_ddr2_memory_pll_sharing_pll_locked,                   --                 .pll_locked
			pll_write_clk_pre_phy_clk => m2_ddr2_memory_pll_sharing_pll_write_clk_pre_phy_clk,    --                 .pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk          => m2_ddr2_memory_pll_sharing_pll_addr_cmd_clk,             --                 .pll_addr_cmd_clk
			pll_avl_clk               => m2_ddr2_memory_pll_sharing_pll_avl_clk,                  --                 .pll_avl_clk
			pll_config_clk            => m2_ddr2_memory_pll_sharing_pll_config_clk,               --                 .pll_config_clk
			dll_pll_locked            => m2_ddr2_memory_dll_sharing_dll_pll_locked,               --      dll_sharing.dll_pll_locked
			dll_delayctrl             => m2_ddr2_memory_dll_sharing_dll_delayctrl                 --                 .dll_delayctrl
		);

	nios2_gen2_0 : component MebX_Qsys_Project_nios2_gen2_0
		port map (
			clk                                 => m2_ddr2_memory_afi_half_clk_clk,                            --                       clk.clk
			reset_n                             => rst_controller_012_reset_out_reset_ports_inv,               --                     reset.reset_n
			reset_req                           => rst_controller_012_reset_out_reset_req,                     --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			i_burstcount                        => nios2_gen2_0_instruction_master_burstcount,                 --                          .burstcount
			i_readdatavalid                     => nios2_gen2_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                       --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory : component MebX_Qsys_Project_onchip_memory
		port map (
			clk        => m2_ddr2_memory_afi_half_clk_clk,               --   clk1.clk
			address    => mm_interconnect_1_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_1_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_1_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_1_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_1_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_1_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_1_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_008_reset_out_reset,            -- reset1.reset
			reset_req  => rst_controller_008_reset_out_reset_req,        --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	pio_button : component MebX_Qsys_Project_pio_BUTTON
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_009_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_pio_button_s1_address,      --                  s1.address
			readdata => mm_interconnect_2_pio_button_s1_readdata,     --                    .readdata
			in_port  => button_export                                 -- external_connection.export
		);

	pio_dip : component MebX_Qsys_Project_pio_DIP
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_009_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_pio_dip_s1_address,         --                  s1.address
			readdata => mm_interconnect_2_pio_dip_s1_readdata,        --                    .readdata
			in_port  => dip_export                                    -- external_connection.export
		);

	pio_ext : component MebX_Qsys_Project_pio_EXT
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_009_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_pio_ext_s1_address,         --                  s1.address
			readdata => mm_interconnect_2_pio_ext_s1_readdata,        --                    .readdata
			in_port  => ext_export                                    -- external_connection.export
		);

	pio_led : component MebX_Qsys_Project_pio_LED
		port map (
			clk        => clk50_clk,                                    --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_2_pio_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_pio_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_pio_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_pio_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_pio_led_s1_readdata,        --                    .readdata
			out_port   => led_de4_export                                -- external_connection.export
		);

	pio_led_painel : component MebX_Qsys_Project_pio_LED_painel
		port map (
			clk        => clk50_clk,                                           --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_2_pio_led_painel_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_pio_led_painel_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_pio_led_painel_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_pio_led_painel_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_pio_led_painel_s1_readdata,        --                    .readdata
			out_port   => led_painel_export                                    -- external_connection.export
		);

	pio_ctrl_io_lvds : component MebX_Qsys_Project_pio_ctrl_io_lvds
		port map (
			clk        => clk50_clk,                                             --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_2_pio_ctrl_io_lvds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_pio_ctrl_io_lvds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_pio_ctrl_io_lvds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_pio_ctrl_io_lvds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_pio_ctrl_io_lvds_s1_readdata,        --                    .readdata
			out_port   => ctrl_io_lvds_export                                    -- external_connection.export
		);

	rmap_mem_nfee_comm_1 : component nrme_rmap_memory_nfee_area_top
		port map (
			reset_i                           => rst_controller_002_reset_out_reset,                                           --                   reset_sink.reset
			clk_100_i                         => m2_ddr2_memory_afi_half_clk_clk,                                              --            clock_sink_100mhz.clk
			avs_0_rmap_address_i              => mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_address,           --          avalon_rmap_slave_0.address
			avs_0_rmap_write_i                => mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_write,             --                             .write
			avs_0_rmap_read_i                 => mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_read,              --                             .read
			avs_0_rmap_readdata_o             => mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_readdata,          --                             .readdata
			avs_0_rmap_writedata_i            => mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_writedata,         --                             .writedata
			avs_0_rmap_waitrequest_o          => mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_waitrequest,       --                             .waitrequest
			avs_0_rmap_byteenable_i           => mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_byteenable,        --                             .byteenable
			fee_0_rmap_wr_address_i           => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_wr_address_signal,    -- conduit_end_fee_rmap_slave_0.wr_address_signal
			fee_0_rmap_write_i                => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_write_signal,         --                             .write_signal
			fee_0_rmap_writedata_i            => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_writedata_signal,     --                             .writedata_signal
			fee_0_rmap_rd_address_i           => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_rd_address_signal,    --                             .rd_address_signal
			fee_0_rmap_read_i                 => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_codec_read_signal,          --                             .read_signal
			fee_0_rmap_wr_waitrequest_o       => rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal,      --                             .wr_waitrequest_signal
			fee_0_rmap_readdata_o             => rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_readdata_signal,            --                             .readdata_signal
			fee_0_rmap_rd_waitrequest_o       => rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal,      --                             .rd_waitrequest_signal
			fee_1_rmap_wr_address_i           => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_wr_address_signal,       -- conduit_end_fee_rmap_slave_1.wr_address_signal
			fee_1_rmap_write_i                => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_write_signal,            --                             .write_signal
			fee_1_rmap_writedata_i            => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_writedata_signal,        --                             .writedata_signal
			fee_1_rmap_rd_address_i           => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_rd_address_signal,       --                             .rd_address_signal
			fee_1_rmap_read_i                 => comm_pedreiro_v1_01_a_conduit_end_fee_rmap_master_hk_read_signal,             --                             .read_signal
			fee_1_rmap_wr_waitrequest_o       => rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal,      --                             .wr_waitrequest_signal
			fee_1_rmap_readdata_o             => rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_readdata_signal,            --                             .readdata_signal
			fee_1_rmap_rd_waitrequest_o       => rmap_mem_nfee_comm_1_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal,      --                             .rd_waitrequest_signal
			channel_hk_timecode_control_i     => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_timecode_control_signal,     --    conduit_end_channel_hk_in.timecode_control_signal
			channel_hk_timecode_time_i        => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_timecode_time_signal,        --                             .timecode_time_signal
			channel_hk_rmap_target_status_i   => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_rmap_target_status_signal,   --                             .rmap_target_status_signal
			channel_hk_rmap_target_indicate_i => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_rmap_target_indicate_signal, --                             .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_i  => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_escape_err_signal,  --                             .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_i  => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_credit_err_signal,  --                             .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_i  => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_parity_err_signal,  --                             .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_i  => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_disconnect_signal,  --                             .spw_link_disconnect_signal
			channel_hk_spw_link_running_i     => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_spw_link_running_signal,     --                             .spw_link_running_signal
			channel_hk_frame_counter_i        => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_frame_counter_signal,        --                             .frame_counter_signal
			channel_hk_frame_number_i         => comm_pedreiro_v1_01_a_conduit_end_channel_hk_out_frame_number_signal,         --                             .frame_number_signal
			avm_rmap_readdata_i               => rmap_mem_nfee_comm_1_avalon_mm_rmap_master_readdata,                          --        avalon_mm_rmap_master.readdata
			avm_rmap_waitrequest_i            => rmap_mem_nfee_comm_1_avalon_mm_rmap_master_waitrequest,                       --                             .waitrequest
			avm_rmap_address_o                => rmap_mem_nfee_comm_1_avalon_mm_rmap_master_address,                           --                             .address
			avm_rmap_read_o                   => rmap_mem_nfee_comm_1_avalon_mm_rmap_master_read,                              --                             .read
			avm_rmap_write_o                  => rmap_mem_nfee_comm_1_avalon_mm_rmap_master_write,                             --                             .write
			avm_rmap_writedata_o              => rmap_mem_nfee_comm_1_avalon_mm_rmap_master_writedata,                         --                             .writedata
			channel_win_mem_addr_offset_i     => comm_pedreiro_v1_01_a_conduit_end_avm_configs_out_win_mem_addr_offset_signal  --   conduit_end_avm_configs_in.win_mem_addr_offset_signal
		);

	rmap_mem_nfee_comm_2 : component nrme_rmap_memory_nfee_area_top
		port map (
			reset_i                           => rst_controller_003_reset_out_reset,                                           --                   reset_sink.reset
			clk_100_i                         => m2_ddr2_memory_afi_half_clk_clk,                                              --            clock_sink_100mhz.clk
			avs_0_rmap_address_i              => mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_address,           --          avalon_rmap_slave_0.address
			avs_0_rmap_write_i                => mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_write,             --                             .write
			avs_0_rmap_read_i                 => mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_read,              --                             .read
			avs_0_rmap_readdata_o             => mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_readdata,          --                             .readdata
			avs_0_rmap_writedata_i            => mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_writedata,         --                             .writedata
			avs_0_rmap_waitrequest_o          => mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_waitrequest,       --                             .waitrequest
			avs_0_rmap_byteenable_i           => mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_byteenable,        --                             .byteenable
			fee_0_rmap_wr_address_i           => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_wr_address_signal,    -- conduit_end_fee_rmap_slave_0.wr_address_signal
			fee_0_rmap_write_i                => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_write_signal,         --                             .write_signal
			fee_0_rmap_writedata_i            => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_writedata_signal,     --                             .writedata_signal
			fee_0_rmap_rd_address_i           => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_rd_address_signal,    --                             .rd_address_signal
			fee_0_rmap_read_i                 => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_codec_read_signal,          --                             .read_signal
			fee_0_rmap_wr_waitrequest_o       => rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal,      --                             .wr_waitrequest_signal
			fee_0_rmap_readdata_o             => rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_readdata_signal,            --                             .readdata_signal
			fee_0_rmap_rd_waitrequest_o       => rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal,      --                             .rd_waitrequest_signal
			fee_1_rmap_wr_address_i           => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_wr_address_signal,       -- conduit_end_fee_rmap_slave_1.wr_address_signal
			fee_1_rmap_write_i                => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_write_signal,            --                             .write_signal
			fee_1_rmap_writedata_i            => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_writedata_signal,        --                             .writedata_signal
			fee_1_rmap_rd_address_i           => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_rd_address_signal,       --                             .rd_address_signal
			fee_1_rmap_read_i                 => comm_pedreiro_v1_01_b_conduit_end_fee_rmap_master_hk_read_signal,             --                             .read_signal
			fee_1_rmap_wr_waitrequest_o       => rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal,      --                             .wr_waitrequest_signal
			fee_1_rmap_readdata_o             => rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_readdata_signal,            --                             .readdata_signal
			fee_1_rmap_rd_waitrequest_o       => rmap_mem_nfee_comm_2_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal,      --                             .rd_waitrequest_signal
			channel_hk_timecode_control_i     => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_timecode_control_signal,     --    conduit_end_channel_hk_in.timecode_control_signal
			channel_hk_timecode_time_i        => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_timecode_time_signal,        --                             .timecode_time_signal
			channel_hk_rmap_target_status_i   => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_rmap_target_status_signal,   --                             .rmap_target_status_signal
			channel_hk_rmap_target_indicate_i => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_rmap_target_indicate_signal, --                             .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_i  => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_escape_err_signal,  --                             .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_i  => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_credit_err_signal,  --                             .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_i  => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_parity_err_signal,  --                             .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_i  => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_disconnect_signal,  --                             .spw_link_disconnect_signal
			channel_hk_spw_link_running_i     => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_spw_link_running_signal,     --                             .spw_link_running_signal
			channel_hk_frame_counter_i        => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_frame_counter_signal,        --                             .frame_counter_signal
			channel_hk_frame_number_i         => comm_pedreiro_v1_01_b_conduit_end_channel_hk_out_frame_number_signal,         --                             .frame_number_signal
			avm_rmap_readdata_i               => rmap_mem_nfee_comm_2_avalon_mm_rmap_master_readdata,                          --        avalon_mm_rmap_master.readdata
			avm_rmap_waitrequest_i            => rmap_mem_nfee_comm_2_avalon_mm_rmap_master_waitrequest,                       --                             .waitrequest
			avm_rmap_address_o                => rmap_mem_nfee_comm_2_avalon_mm_rmap_master_address,                           --                             .address
			avm_rmap_read_o                   => rmap_mem_nfee_comm_2_avalon_mm_rmap_master_read,                              --                             .read
			avm_rmap_write_o                  => rmap_mem_nfee_comm_2_avalon_mm_rmap_master_write,                             --                             .write
			avm_rmap_writedata_o              => rmap_mem_nfee_comm_2_avalon_mm_rmap_master_writedata,                         --                             .writedata
			channel_win_mem_addr_offset_i     => comm_pedreiro_v1_01_b_conduit_end_avm_configs_out_win_mem_addr_offset_signal  --   conduit_end_avm_configs_in.win_mem_addr_offset_signal
		);

	rmap_mem_nfee_comm_3 : component nrme_rmap_memory_nfee_area_top
		port map (
			reset_i                           => rst_controller_004_reset_out_reset,                                           --                   reset_sink.reset
			clk_100_i                         => m2_ddr2_memory_afi_half_clk_clk,                                              --            clock_sink_100mhz.clk
			avs_0_rmap_address_i              => mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_address,           --          avalon_rmap_slave_0.address
			avs_0_rmap_write_i                => mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_write,             --                             .write
			avs_0_rmap_read_i                 => mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_read,              --                             .read
			avs_0_rmap_readdata_o             => mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_readdata,          --                             .readdata
			avs_0_rmap_writedata_i            => mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_writedata,         --                             .writedata
			avs_0_rmap_waitrequest_o          => mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_waitrequest,       --                             .waitrequest
			avs_0_rmap_byteenable_i           => mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_byteenable,        --                             .byteenable
			fee_0_rmap_wr_address_i           => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_wr_address_signal,    -- conduit_end_fee_rmap_slave_0.wr_address_signal
			fee_0_rmap_write_i                => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_write_signal,         --                             .write_signal
			fee_0_rmap_writedata_i            => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_writedata_signal,     --                             .writedata_signal
			fee_0_rmap_rd_address_i           => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_rd_address_signal,    --                             .rd_address_signal
			fee_0_rmap_read_i                 => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_codec_read_signal,          --                             .read_signal
			fee_0_rmap_wr_waitrequest_o       => rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal,      --                             .wr_waitrequest_signal
			fee_0_rmap_readdata_o             => rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_readdata_signal,            --                             .readdata_signal
			fee_0_rmap_rd_waitrequest_o       => rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal,      --                             .rd_waitrequest_signal
			fee_1_rmap_wr_address_i           => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_wr_address_signal,       -- conduit_end_fee_rmap_slave_1.wr_address_signal
			fee_1_rmap_write_i                => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_write_signal,            --                             .write_signal
			fee_1_rmap_writedata_i            => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_writedata_signal,        --                             .writedata_signal
			fee_1_rmap_rd_address_i           => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_rd_address_signal,       --                             .rd_address_signal
			fee_1_rmap_read_i                 => comm_pedreiro_v1_01_c_conduit_end_fee_rmap_master_hk_read_signal,             --                             .read_signal
			fee_1_rmap_wr_waitrequest_o       => rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal,      --                             .wr_waitrequest_signal
			fee_1_rmap_readdata_o             => rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_readdata_signal,            --                             .readdata_signal
			fee_1_rmap_rd_waitrequest_o       => rmap_mem_nfee_comm_3_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal,      --                             .rd_waitrequest_signal
			channel_hk_timecode_control_i     => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_timecode_control_signal,     --    conduit_end_channel_hk_in.timecode_control_signal
			channel_hk_timecode_time_i        => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_timecode_time_signal,        --                             .timecode_time_signal
			channel_hk_rmap_target_status_i   => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_rmap_target_status_signal,   --                             .rmap_target_status_signal
			channel_hk_rmap_target_indicate_i => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_rmap_target_indicate_signal, --                             .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_i  => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_escape_err_signal,  --                             .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_i  => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_credit_err_signal,  --                             .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_i  => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_parity_err_signal,  --                             .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_i  => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_disconnect_signal,  --                             .spw_link_disconnect_signal
			channel_hk_spw_link_running_i     => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_spw_link_running_signal,     --                             .spw_link_running_signal
			channel_hk_frame_counter_i        => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_frame_counter_signal,        --                             .frame_counter_signal
			channel_hk_frame_number_i         => comm_pedreiro_v1_01_c_conduit_end_channel_hk_out_frame_number_signal,         --                             .frame_number_signal
			avm_rmap_readdata_i               => rmap_mem_nfee_comm_3_avalon_mm_rmap_master_readdata,                          --        avalon_mm_rmap_master.readdata
			avm_rmap_waitrequest_i            => rmap_mem_nfee_comm_3_avalon_mm_rmap_master_waitrequest,                       --                             .waitrequest
			avm_rmap_address_o                => rmap_mem_nfee_comm_3_avalon_mm_rmap_master_address,                           --                             .address
			avm_rmap_read_o                   => rmap_mem_nfee_comm_3_avalon_mm_rmap_master_read,                              --                             .read
			avm_rmap_write_o                  => rmap_mem_nfee_comm_3_avalon_mm_rmap_master_write,                             --                             .write
			avm_rmap_writedata_o              => rmap_mem_nfee_comm_3_avalon_mm_rmap_master_writedata,                         --                             .writedata
			channel_win_mem_addr_offset_i     => comm_pedreiro_v1_01_c_conduit_end_avm_configs_out_win_mem_addr_offset_signal  --   conduit_end_avm_configs_in.win_mem_addr_offset_signal
		);

	rmap_mem_nfee_comm_4 : component nrme_rmap_memory_nfee_area_top
		port map (
			reset_i                           => rst_controller_005_reset_out_reset,                                           --                   reset_sink.reset
			clk_100_i                         => m2_ddr2_memory_afi_half_clk_clk,                                              --            clock_sink_100mhz.clk
			avs_0_rmap_address_i              => mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_address,           --          avalon_rmap_slave_0.address
			avs_0_rmap_write_i                => mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_write,             --                             .write
			avs_0_rmap_read_i                 => mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_read,              --                             .read
			avs_0_rmap_readdata_o             => mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_readdata,          --                             .readdata
			avs_0_rmap_writedata_i            => mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_writedata,         --                             .writedata
			avs_0_rmap_waitrequest_o          => mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_waitrequest,       --                             .waitrequest
			avs_0_rmap_byteenable_i           => mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_byteenable,        --                             .byteenable
			fee_0_rmap_wr_address_i           => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_wr_address_signal,    -- conduit_end_fee_rmap_slave_0.wr_address_signal
			fee_0_rmap_write_i                => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_write_signal,         --                             .write_signal
			fee_0_rmap_writedata_i            => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_writedata_signal,     --                             .writedata_signal
			fee_0_rmap_rd_address_i           => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_rd_address_signal,    --                             .rd_address_signal
			fee_0_rmap_read_i                 => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_codec_read_signal,          --                             .read_signal
			fee_0_rmap_wr_waitrequest_o       => rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal,      --                             .wr_waitrequest_signal
			fee_0_rmap_readdata_o             => rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_readdata_signal,            --                             .readdata_signal
			fee_0_rmap_rd_waitrequest_o       => rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal,      --                             .rd_waitrequest_signal
			fee_1_rmap_wr_address_i           => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_wr_address_signal,       -- conduit_end_fee_rmap_slave_1.wr_address_signal
			fee_1_rmap_write_i                => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_write_signal,            --                             .write_signal
			fee_1_rmap_writedata_i            => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_writedata_signal,        --                             .writedata_signal
			fee_1_rmap_rd_address_i           => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_rd_address_signal,       --                             .rd_address_signal
			fee_1_rmap_read_i                 => comm_pedreiro_v1_01_d_conduit_end_fee_rmap_master_hk_read_signal,             --                             .read_signal
			fee_1_rmap_wr_waitrequest_o       => rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal,      --                             .wr_waitrequest_signal
			fee_1_rmap_readdata_o             => rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_readdata_signal,            --                             .readdata_signal
			fee_1_rmap_rd_waitrequest_o       => rmap_mem_nfee_comm_4_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal,      --                             .rd_waitrequest_signal
			channel_hk_timecode_control_i     => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_timecode_control_signal,     --    conduit_end_channel_hk_in.timecode_control_signal
			channel_hk_timecode_time_i        => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_timecode_time_signal,        --                             .timecode_time_signal
			channel_hk_rmap_target_status_i   => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_rmap_target_status_signal,   --                             .rmap_target_status_signal
			channel_hk_rmap_target_indicate_i => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_rmap_target_indicate_signal, --                             .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_i  => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_escape_err_signal,  --                             .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_i  => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_credit_err_signal,  --                             .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_i  => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_parity_err_signal,  --                             .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_i  => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_disconnect_signal,  --                             .spw_link_disconnect_signal
			channel_hk_spw_link_running_i     => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_spw_link_running_signal,     --                             .spw_link_running_signal
			channel_hk_frame_counter_i        => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_frame_counter_signal,        --                             .frame_counter_signal
			channel_hk_frame_number_i         => comm_pedreiro_v1_01_d_conduit_end_channel_hk_out_frame_number_signal,         --                             .frame_number_signal
			avm_rmap_readdata_i               => rmap_mem_nfee_comm_4_avalon_mm_rmap_master_readdata,                          --        avalon_mm_rmap_master.readdata
			avm_rmap_waitrequest_i            => rmap_mem_nfee_comm_4_avalon_mm_rmap_master_waitrequest,                       --                             .waitrequest
			avm_rmap_address_o                => rmap_mem_nfee_comm_4_avalon_mm_rmap_master_address,                           --                             .address
			avm_rmap_read_o                   => rmap_mem_nfee_comm_4_avalon_mm_rmap_master_read,                              --                             .read
			avm_rmap_write_o                  => rmap_mem_nfee_comm_4_avalon_mm_rmap_master_write,                             --                             .write
			avm_rmap_writedata_o              => rmap_mem_nfee_comm_4_avalon_mm_rmap_master_writedata,                         --                             .writedata
			channel_win_mem_addr_offset_i     => comm_pedreiro_v1_01_d_conduit_end_avm_configs_out_win_mem_addr_offset_signal  --   conduit_end_avm_configs_in.win_mem_addr_offset_signal
		);

	rmap_mem_nfee_comm_5 : component nrme_rmap_memory_nfee_area_top
		port map (
			reset_i                           => rst_controller_006_reset_out_reset,                                           --                   reset_sink.reset
			clk_100_i                         => m2_ddr2_memory_afi_half_clk_clk,                                              --            clock_sink_100mhz.clk
			avs_0_rmap_address_i              => mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_address,           --          avalon_rmap_slave_0.address
			avs_0_rmap_write_i                => mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_write,             --                             .write
			avs_0_rmap_read_i                 => mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_read,              --                             .read
			avs_0_rmap_readdata_o             => mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_readdata,          --                             .readdata
			avs_0_rmap_writedata_i            => mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_writedata,         --                             .writedata
			avs_0_rmap_waitrequest_o          => mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_waitrequest,       --                             .waitrequest
			avs_0_rmap_byteenable_i           => mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_byteenable,        --                             .byteenable
			fee_0_rmap_wr_address_i           => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_wr_address_signal,    -- conduit_end_fee_rmap_slave_0.wr_address_signal
			fee_0_rmap_write_i                => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_write_signal,         --                             .write_signal
			fee_0_rmap_writedata_i            => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_writedata_signal,     --                             .writedata_signal
			fee_0_rmap_rd_address_i           => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_rd_address_signal,    --                             .rd_address_signal
			fee_0_rmap_read_i                 => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_codec_read_signal,          --                             .read_signal
			fee_0_rmap_wr_waitrequest_o       => rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal,      --                             .wr_waitrequest_signal
			fee_0_rmap_readdata_o             => rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_readdata_signal,            --                             .readdata_signal
			fee_0_rmap_rd_waitrequest_o       => rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal,      --                             .rd_waitrequest_signal
			fee_1_rmap_wr_address_i           => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_wr_address_signal,       -- conduit_end_fee_rmap_slave_1.wr_address_signal
			fee_1_rmap_write_i                => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_write_signal,            --                             .write_signal
			fee_1_rmap_writedata_i            => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_writedata_signal,        --                             .writedata_signal
			fee_1_rmap_rd_address_i           => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_rd_address_signal,       --                             .rd_address_signal
			fee_1_rmap_read_i                 => comm_pedreiro_v1_01_e_conduit_end_fee_rmap_master_hk_read_signal,             --                             .read_signal
			fee_1_rmap_wr_waitrequest_o       => rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal,      --                             .wr_waitrequest_signal
			fee_1_rmap_readdata_o             => rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_readdata_signal,            --                             .readdata_signal
			fee_1_rmap_rd_waitrequest_o       => rmap_mem_nfee_comm_5_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal,      --                             .rd_waitrequest_signal
			channel_hk_timecode_control_i     => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_timecode_control_signal,     --    conduit_end_channel_hk_in.timecode_control_signal
			channel_hk_timecode_time_i        => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_timecode_time_signal,        --                             .timecode_time_signal
			channel_hk_rmap_target_status_i   => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_rmap_target_status_signal,   --                             .rmap_target_status_signal
			channel_hk_rmap_target_indicate_i => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_rmap_target_indicate_signal, --                             .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_i  => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_escape_err_signal,  --                             .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_i  => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_credit_err_signal,  --                             .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_i  => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_parity_err_signal,  --                             .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_i  => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_disconnect_signal,  --                             .spw_link_disconnect_signal
			channel_hk_spw_link_running_i     => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_spw_link_running_signal,     --                             .spw_link_running_signal
			channel_hk_frame_counter_i        => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_frame_counter_signal,        --                             .frame_counter_signal
			channel_hk_frame_number_i         => comm_pedreiro_v1_01_e_conduit_end_channel_hk_out_frame_number_signal,         --                             .frame_number_signal
			avm_rmap_readdata_i               => rmap_mem_nfee_comm_5_avalon_mm_rmap_master_readdata,                          --        avalon_mm_rmap_master.readdata
			avm_rmap_waitrequest_i            => rmap_mem_nfee_comm_5_avalon_mm_rmap_master_waitrequest,                       --                             .waitrequest
			avm_rmap_address_o                => rmap_mem_nfee_comm_5_avalon_mm_rmap_master_address,                           --                             .address
			avm_rmap_read_o                   => rmap_mem_nfee_comm_5_avalon_mm_rmap_master_read,                              --                             .read
			avm_rmap_write_o                  => rmap_mem_nfee_comm_5_avalon_mm_rmap_master_write,                             --                             .write
			avm_rmap_writedata_o              => rmap_mem_nfee_comm_5_avalon_mm_rmap_master_writedata,                         --                             .writedata
			channel_win_mem_addr_offset_i     => comm_pedreiro_v1_01_e_conduit_end_avm_configs_out_win_mem_addr_offset_signal  --   conduit_end_avm_configs_in.win_mem_addr_offset_signal
		);

	rmap_mem_nfee_comm_6 : component nrme_rmap_memory_nfee_area_top
		port map (
			reset_i                           => rst_controller_007_reset_out_reset,                                           --                   reset_sink.reset
			clk_100_i                         => m2_ddr2_memory_afi_half_clk_clk,                                              --            clock_sink_100mhz.clk
			avs_0_rmap_address_i              => mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_address,           --          avalon_rmap_slave_0.address
			avs_0_rmap_write_i                => mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_write,             --                             .write
			avs_0_rmap_read_i                 => mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_read,              --                             .read
			avs_0_rmap_readdata_o             => mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_readdata,          --                             .readdata
			avs_0_rmap_writedata_i            => mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_writedata,         --                             .writedata
			avs_0_rmap_waitrequest_o          => mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_waitrequest,       --                             .waitrequest
			avs_0_rmap_byteenable_i           => mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_byteenable,        --                             .byteenable
			fee_0_rmap_wr_address_i           => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_wr_address_signal,    -- conduit_end_fee_rmap_slave_0.wr_address_signal
			fee_0_rmap_write_i                => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_write_signal,         --                             .write_signal
			fee_0_rmap_writedata_i            => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_writedata_signal,     --                             .writedata_signal
			fee_0_rmap_rd_address_i           => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_rd_address_signal,    --                             .rd_address_signal
			fee_0_rmap_read_i                 => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_codec_read_signal,          --                             .read_signal
			fee_0_rmap_wr_waitrequest_o       => rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_wr_waitrequest_signal,      --                             .wr_waitrequest_signal
			fee_0_rmap_readdata_o             => rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_readdata_signal,            --                             .readdata_signal
			fee_0_rmap_rd_waitrequest_o       => rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_0_rd_waitrequest_signal,      --                             .rd_waitrequest_signal
			fee_1_rmap_wr_address_i           => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_wr_address_signal,       -- conduit_end_fee_rmap_slave_1.wr_address_signal
			fee_1_rmap_write_i                => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_write_signal,            --                             .write_signal
			fee_1_rmap_writedata_i            => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_writedata_signal,        --                             .writedata_signal
			fee_1_rmap_rd_address_i           => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_rd_address_signal,       --                             .rd_address_signal
			fee_1_rmap_read_i                 => comm_pedreiro_v1_01_f_conduit_end_fee_rmap_master_hk_read_signal,             --                             .read_signal
			fee_1_rmap_wr_waitrequest_o       => rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_wr_waitrequest_signal,      --                             .wr_waitrequest_signal
			fee_1_rmap_readdata_o             => rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_readdata_signal,            --                             .readdata_signal
			fee_1_rmap_rd_waitrequest_o       => rmap_mem_nfee_comm_6_conduit_end_fee_rmap_slave_1_rd_waitrequest_signal,      --                             .rd_waitrequest_signal
			channel_hk_timecode_control_i     => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_timecode_control_signal,     --    conduit_end_channel_hk_in.timecode_control_signal
			channel_hk_timecode_time_i        => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_timecode_time_signal,        --                             .timecode_time_signal
			channel_hk_rmap_target_status_i   => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_rmap_target_status_signal,   --                             .rmap_target_status_signal
			channel_hk_rmap_target_indicate_i => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_rmap_target_indicate_signal, --                             .rmap_target_indicate_signal
			channel_hk_spw_link_escape_err_i  => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_escape_err_signal,  --                             .spw_link_escape_err_signal
			channel_hk_spw_link_credit_err_i  => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_credit_err_signal,  --                             .spw_link_credit_err_signal
			channel_hk_spw_link_parity_err_i  => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_parity_err_signal,  --                             .spw_link_parity_err_signal
			channel_hk_spw_link_disconnect_i  => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_disconnect_signal,  --                             .spw_link_disconnect_signal
			channel_hk_spw_link_running_i     => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_spw_link_running_signal,     --                             .spw_link_running_signal
			channel_hk_frame_counter_i        => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_frame_counter_signal,        --                             .frame_counter_signal
			channel_hk_frame_number_i         => comm_pedreiro_v1_01_f_conduit_end_channel_hk_out_frame_number_signal,         --                             .frame_number_signal
			avm_rmap_readdata_i               => rmap_mem_nfee_comm_6_avalon_mm_rmap_master_readdata,                          --        avalon_mm_rmap_master.readdata
			avm_rmap_waitrequest_i            => rmap_mem_nfee_comm_6_avalon_mm_rmap_master_waitrequest,                       --                             .waitrequest
			avm_rmap_address_o                => rmap_mem_nfee_comm_6_avalon_mm_rmap_master_address,                           --                             .address
			avm_rmap_read_o                   => rmap_mem_nfee_comm_6_avalon_mm_rmap_master_read,                              --                             .read
			avm_rmap_write_o                  => rmap_mem_nfee_comm_6_avalon_mm_rmap_master_write,                             --                             .write
			avm_rmap_writedata_o              => rmap_mem_nfee_comm_6_avalon_mm_rmap_master_writedata,                         --                             .writedata
			channel_win_mem_addr_offset_i     => comm_pedreiro_v1_01_f_conduit_end_avm_configs_out_win_mem_addr_offset_signal  --   conduit_end_avm_configs_in.win_mem_addr_offset_signal
		);

	rs232_uart : component MebX_Qsys_Project_rs232_uart
		port map (
			clk           => clk50_clk,                                       --                 clk.clk
			reset_n       => rst_controller_013_reset_out_reset_ports_inv,    --               reset.reset_n
			address       => mm_interconnect_2_rs232_uart_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_2_rs232_uart_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_2_rs232_uart_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_2_rs232_uart_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_2_rs232_uart_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_2_rs232_uart_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_2_rs232_uart_s1_readdata,        --                    .readdata
			rxd           => rs232_uart_rxd,                                  -- external_connection.export
			txd           => rs232_uart_txd,                                  --                    .export
			irq           => irq_synchronizer_002_receiver_irq(0)             --                 irq.irq
		);

	rst_controller : component rst_controller_top
		port map (
			clock_sink_clk                          => clk50_clk,                                                                --                  clock_sink.clk
			reset_sink_reset                        => rst_controller_009_reset_out_reset,                                       --                  reset_sink.reset
			reset_source_ftdi_reset                 => open,                                                                     --           reset_source_ftdi.reset
			reset_source_sync_reset                 => rst_controller_reset_source_sync_reset,                                   --           reset_source_sync.reset
			reset_source_rs232_reset                => rst_controller_reset_source_rs232_reset,                                  --          reset_source_rs232.reset
			reset_source_sd_card_reset              => rst_controller_reset_source_sd_card_reset,                                --        reset_source_sd_card.reset
			reset_source_comm_ch8_reset             => open,                                                                     --       reset_source_comm_ch8.reset
			reset_source_comm_ch7_reset             => open,                                                                     --       reset_source_comm_ch7.reset
			reset_source_comm_ch6_reset             => rst_controller_reset_source_comm_ch6_reset,                               --       reset_source_comm_ch6.reset
			reset_source_comm_ch5_reset             => rst_controller_reset_source_comm_ch5_reset,                               --       reset_source_comm_ch5.reset
			reset_source_comm_ch4_reset             => rst_controller_reset_source_comm_ch4_reset,                               --       reset_source_comm_ch4.reset
			reset_source_comm_ch3_reset             => rst_controller_reset_source_comm_ch3_reset,                               --       reset_source_comm_ch3.reset
			reset_source_comm_ch2_reset             => rst_controller_reset_source_comm_ch2_reset,                               --       reset_source_comm_ch2.reset
			reset_source_comm_ch1_reset             => rst_controller_reset_source_comm_ch1_reset,                               --       reset_source_comm_ch1.reset
			avalon_slave_rst_controller_address     => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_address,     -- avalon_rst_controller_slave.address
			avalon_slave_rst_controller_write       => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_write,       --                            .write
			avalon_slave_rst_controller_read        => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_read,        --                            .read
			avalon_slave_rst_controller_writedata   => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_writedata,   --                            .writedata
			avalon_slave_rst_controller_readdata    => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_readdata,    --                            .readdata
			avalon_slave_rst_controller_waitrequest => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_waitrequest, --                            .waitrequest
			simucam_reset_signal                    => rst_controller_conduit_simucam_reset_t_simucam_reset_signal,              --       conduit_simucam_reset.t_simucam_reset_signal
			reset_input_signal                      => rst_controller_conduit_reset_input_t_reset_input_signal                   --         conduit_reset_input.t_reset_input_signal
		);

	rtcc_alarm : component MebX_Qsys_Project_csense_sdo
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_009_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_rtcc_alarm_s1_address,      --                  s1.address
			readdata => mm_interconnect_2_rtcc_alarm_s1_readdata,     --                    .readdata
			in_port  => rtcc_alarm_export                             -- external_connection.export
		);

	rtcc_cs_n : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                      --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_2_rtcc_cs_n_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_rtcc_cs_n_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_rtcc_cs_n_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_rtcc_cs_n_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_rtcc_cs_n_s1_readdata,        --                    .readdata
			out_port   => rtcc_cs_n_export                                -- external_connection.export
		);

	rtcc_sck : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                     --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_2_rtcc_sck_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_rtcc_sck_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_rtcc_sck_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_rtcc_sck_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_rtcc_sck_s1_readdata,        --                    .readdata
			out_port   => rtcc_sck_export                                -- external_connection.export
		);

	rtcc_sdi : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                     --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_2_rtcc_sdi_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_rtcc_sdi_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_rtcc_sdi_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_rtcc_sdi_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_rtcc_sdi_s1_readdata,        --                    .readdata
			out_port   => rtcc_sdi_export                                -- external_connection.export
		);

	rtcc_sdo : component MebX_Qsys_Project_csense_sdo
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_009_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_rtcc_sdo_s1_address,        --                  s1.address
			readdata => mm_interconnect_2_rtcc_sdo_s1_readdata,       --                    .readdata
			in_port  => rtcc_sdo_export                               -- external_connection.export
		);

	sd_card_wp_n : component MebX_Qsys_Project_csense_sdo
		port map (
			clk      => clk50_clk,                                    --                 clk.clk
			reset_n  => rst_controller_009_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_2_sd_card_wp_n_s1_address,    --                  s1.address
			readdata => mm_interconnect_2_sd_card_wp_n_s1_readdata,   --                    .readdata
			in_port  => sd_card_wp_n_io_export                        -- external_connection.export
		);

	sync : component sync_ent
		generic map (
			g_SYNC_IRQ_NUMBER     => 11,
			g_PRE_SYNC_IRQ_NUMBER => 12
		)
		port map (
			clock_sink_clk_i                => clk50_clk,                                          --                     clock.clk
			reset_sink_reset_i              => rst_controller_014_reset_out_reset,                 --                     reset.reset
			avalon_slave_address_i          => mm_interconnect_2_sync_avalon_mm_slave_address,     --           avalon_mm_slave.address
			avalon_slave_read_i             => mm_interconnect_2_sync_avalon_mm_slave_read,        --                          .read
			avalon_slave_write_i            => mm_interconnect_2_sync_avalon_mm_slave_write,       --                          .write
			avalon_slave_writedata_i        => mm_interconnect_2_sync_avalon_mm_slave_writedata,   --                          .writedata
			avalon_slave_byteenable_i       => mm_interconnect_2_sync_avalon_mm_slave_byteenable,  --                          .byteenable
			avalon_slave_readdata_o         => mm_interconnect_2_sync_avalon_mm_slave_readdata,    --                          .readdata
			avalon_slave_waitrequest_o      => mm_interconnect_2_sync_avalon_mm_slave_waitrequest, --                          .waitrequest
			conduit_sync_signal_syncin_i    => sync_in_conduit,                                    --                   sync_in.conduit
			conduit_sync_signal_spw1_o      => sync_spw1_conduit,                                  --                 sync_spw1.conduit
			conduit_sync_signal_spw2_o      => sync_spw2_conduit,                                  --                 sync_spw2.conduit
			conduit_sync_signal_spw3_o      => sync_spw3_conduit,                                  --                 sync_spw3.conduit
			conduit_sync_signal_spw4_o      => sync_spw4_conduit,                                  --                 sync_spw4.conduit
			conduit_sync_signal_spw5_o      => sync_spw5_conduit,                                  --                 sync_spw5.conduit
			conduit_sync_signal_spw6_o      => sync_spw6_conduit,                                  --                 sync_spw6.conduit
			conduit_sync_signal_spw7_o      => sync_spw7_conduit,                                  --                 sync_spw7.conduit
			conduit_sync_signal_spw8_o      => sync_spw8_conduit,                                  --                 sync_spw8.conduit
			conduit_sync_signal_syncout_o   => sync_out_conduit,                                   --                  sync_out.conduit
			sync_interrupt_sender_irq_o     => irq_synchronizer_004_receiver_irq(0),               --     sync_interrupt_sender.irq
			pre_sync_interrupt_sender_irq_o => irq_synchronizer_003_receiver_irq(0)                -- pre_sync_interrupt_sender.irq
		);

	sysid_qsys : component MebX_Qsys_Project_sysid_qsys
		port map (
			clock    => m2_ddr2_memory_afi_half_clk_clk,                       --           clk.clk
			reset_n  => rst_controller_008_reset_out_reset_ports_inv,          --         reset.reset_n
			readdata => mm_interconnect_1_sysid_qsys_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_1_sysid_qsys_control_slave_address(0)  --              .address
		);

	temp_scl : component MebX_Qsys_Project_csense_adc_fo
		port map (
			clk        => clk50_clk,                                     --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_2_temp_scl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_temp_scl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_temp_scl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_temp_scl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_temp_scl_s1_readdata,        --                    .readdata
			out_port   => temp_scl_export                                -- external_connection.export
		);

	temp_sda : component MebX_Qsys_Project_m1_ddr2_i2c_sda
		port map (
			clk        => clk50_clk,                                     --                 clk.clk
			reset_n    => rst_controller_009_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_2_temp_sda_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_temp_sda_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_temp_sda_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_temp_sda_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_temp_sda_s1_readdata,        --                    .readdata
			bidir_port => temp_sda_export                                -- external_connection.export
		);

	timer_1ms : component MebX_Qsys_Project_timer_1ms
		port map (
			clk           => clk50_clk,                                      --           clk.clk
			reset_n       => rst_controller_009_reset_out_reset_ports_inv,   --         reset.reset_n
			address       => mm_interconnect_2_timer_1ms_s1_address,         --            s1.address
			writedata     => mm_interconnect_2_timer_1ms_s1_writedata,       --              .writedata
			readdata      => mm_interconnect_2_timer_1ms_s1_readdata,        --              .readdata
			chipselect    => mm_interconnect_2_timer_1ms_s1_chipselect,      --              .chipselect
			write_n       => mm_interconnect_2_timer_1ms_s1_write_ports_inv, --              .write_n
			irq           => irq_synchronizer_receiver_irq(0),               --           irq.irq
			timeout_pulse => timer_1ms_external_port_export                  -- external_port.export
		);

	timer_1us : component MebX_Qsys_Project_timer_1us
		port map (
			clk           => clk50_clk,                                      --           clk.clk
			reset_n       => rst_controller_009_reset_out_reset_ports_inv,   --         reset.reset_n
			address       => mm_interconnect_2_timer_1us_s1_address,         --            s1.address
			writedata     => mm_interconnect_2_timer_1us_s1_writedata,       --              .writedata
			readdata      => mm_interconnect_2_timer_1us_s1_readdata,        --              .readdata
			chipselect    => mm_interconnect_2_timer_1us_s1_chipselect,      --              .chipselect
			write_n       => mm_interconnect_2_timer_1us_s1_write_ports_inv, --              .write_n
			irq           => irq_synchronizer_001_receiver_irq(0),           --           irq.irq
			timeout_pulse => timer_1us_external_port_export                  -- external_port.export
		);

	tristate_conduit_bridge_0 : component MebX_Qsys_Project_tristate_conduit_bridge_0
		port map (
			clk                         => m2_ddr2_memory_afi_half_clk_clk,       --   clk.clk
			reset                       => rst_controller_010_reset_out_reset,    -- reset.reset
			request                     => ext_flash_tcm_request,                 --   tcs.request
			grant                       => ext_flash_tcm_grant,                   --      .grant
			tcs_tcm_address_out         => ext_flash_tcm_address_out,             --      .address_out
			tcs_tcm_read_n_out(0)       => ext_flash_tcm_read_n_out,              --      .read_n_out
			tcs_tcm_write_n_out(0)      => ext_flash_tcm_write_n_out,             --      .write_n_out
			tcs_tcm_data_out            => ext_flash_tcm_data_out,                --      .data_out
			tcs_tcm_data_outen          => ext_flash_tcm_data_outen,              --      .data_outen
			tcs_tcm_data_in             => ext_flash_tcm_data_in,                 --      .data_in
			tcs_tcm_chipselect_n_out(0) => ext_flash_tcm_chipselect_n_out,        --      .chipselect_n_out
			tcm_address_out             => tristate_conduit_tcm_address_out,      --   out.tcm_address_out
			tcm_read_n_out              => tristate_conduit_tcm_read_n_out,       --      .tcm_read_n_out
			tcm_write_n_out             => tristate_conduit_tcm_write_n_out,      --      .tcm_write_n_out
			tcm_data_out                => tristate_conduit_tcm_data_out,         --      .tcm_data_out
			tcm_chipselect_n_out        => tristate_conduit_tcm_chipselect_n_out  --      .tcm_chipselect_n_out
		);

	mm_interconnect_0 : component MebX_Qsys_Project_mm_interconnect_0
		port map (
			clk_100_clk_clk                                                 => m2_ddr2_memory_afi_half_clk_clk,                          --                                               clk_100_clk.clk
			m2_ddr2_memory_afi_clk_clk                                      => m2_ddr2_memory_afi_clk_clk,                               --                                    m2_ddr2_memory_afi_clk.clk
			m2_ddr2_memory_afi_half_clk_clk                                 => m2_ddr2_memory_afi_half_clk_clk,                          --                               m2_ddr2_memory_afi_half_clk.clk
			ddr2_address_span_extender_reset_reset_bridge_in_reset_reset    => rst_controller_008_reset_out_reset,                       --    ddr2_address_span_extender_reset_reset_bridge_in_reset.reset
			m1_clock_bridge_s0_reset_reset_bridge_in_reset_reset            => rst_controller_008_reset_out_reset,                       --            m1_clock_bridge_s0_reset_reset_bridge_in_reset.reset
			m2_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset => rst_controller_015_reset_out_reset,                       -- m2_ddr2_memory_avl_translator_reset_reset_bridge_in_reset.reset
			m2_ddr2_memory_soft_reset_reset_bridge_in_reset_reset           => rst_controller_015_reset_out_reset,                       --           m2_ddr2_memory_soft_reset_reset_bridge_in_reset.reset
			rmap_mem_nfee_comm_1_reset_sink_reset_bridge_in_reset_reset     => rst_controller_002_reset_out_reset,                       --     rmap_mem_nfee_comm_1_reset_sink_reset_bridge_in_reset.reset
			rmap_mem_nfee_comm_2_reset_sink_reset_bridge_in_reset_reset     => rst_controller_003_reset_out_reset,                       --     rmap_mem_nfee_comm_2_reset_sink_reset_bridge_in_reset.reset
			rmap_mem_nfee_comm_3_reset_sink_reset_bridge_in_reset_reset     => rst_controller_004_reset_out_reset,                       --     rmap_mem_nfee_comm_3_reset_sink_reset_bridge_in_reset.reset
			rmap_mem_nfee_comm_4_reset_sink_reset_bridge_in_reset_reset     => rst_controller_005_reset_out_reset,                       --     rmap_mem_nfee_comm_4_reset_sink_reset_bridge_in_reset.reset
			rmap_mem_nfee_comm_5_reset_sink_reset_bridge_in_reset_reset     => rst_controller_006_reset_out_reset,                       --     rmap_mem_nfee_comm_5_reset_sink_reset_bridge_in_reset.reset
			rmap_mem_nfee_comm_6_reset_sink_reset_bridge_in_reset_reset     => rst_controller_007_reset_out_reset,                       --     rmap_mem_nfee_comm_6_reset_sink_reset_bridge_in_reset.reset
			ddr2_address_span_extender_expanded_master_address              => ddr2_address_span_extender_expanded_master_address,       --                ddr2_address_span_extender_expanded_master.address
			ddr2_address_span_extender_expanded_master_waitrequest          => ddr2_address_span_extender_expanded_master_waitrequest,   --                                                          .waitrequest
			ddr2_address_span_extender_expanded_master_burstcount           => ddr2_address_span_extender_expanded_master_burstcount,    --                                                          .burstcount
			ddr2_address_span_extender_expanded_master_byteenable           => ddr2_address_span_extender_expanded_master_byteenable,    --                                                          .byteenable
			ddr2_address_span_extender_expanded_master_read                 => ddr2_address_span_extender_expanded_master_read,          --                                                          .read
			ddr2_address_span_extender_expanded_master_readdata             => ddr2_address_span_extender_expanded_master_readdata,      --                                                          .readdata
			ddr2_address_span_extender_expanded_master_readdatavalid        => ddr2_address_span_extender_expanded_master_readdatavalid, --                                                          .readdatavalid
			ddr2_address_span_extender_expanded_master_write                => ddr2_address_span_extender_expanded_master_write,         --                                                          .write
			ddr2_address_span_extender_expanded_master_writedata            => ddr2_address_span_extender_expanded_master_writedata,     --                                                          .writedata
			dma_comm_1_left_mm_read_address                                 => dma_comm_1_left_mm_read_address,                          --                                   dma_comm_1_left_mm_read.address
			dma_comm_1_left_mm_read_waitrequest                             => dma_comm_1_left_mm_read_waitrequest,                      --                                                          .waitrequest
			dma_comm_1_left_mm_read_byteenable                              => dma_comm_1_left_mm_read_byteenable,                       --                                                          .byteenable
			dma_comm_1_left_mm_read_read                                    => dma_comm_1_left_mm_read_read,                             --                                                          .read
			dma_comm_1_left_mm_read_readdata                                => dma_comm_1_left_mm_read_readdata,                         --                                                          .readdata
			dma_comm_1_left_mm_read_readdatavalid                           => dma_comm_1_left_mm_read_readdatavalid,                    --                                                          .readdatavalid
			dma_comm_1_right_mm_read_address                                => dma_comm_1_right_mm_read_address,                         --                                  dma_comm_1_right_mm_read.address
			dma_comm_1_right_mm_read_waitrequest                            => dma_comm_1_right_mm_read_waitrequest,                     --                                                          .waitrequest
			dma_comm_1_right_mm_read_byteenable                             => dma_comm_1_right_mm_read_byteenable,                      --                                                          .byteenable
			dma_comm_1_right_mm_read_read                                   => dma_comm_1_right_mm_read_read,                            --                                                          .read
			dma_comm_1_right_mm_read_readdata                               => dma_comm_1_right_mm_read_readdata,                        --                                                          .readdata
			dma_comm_1_right_mm_read_readdatavalid                          => dma_comm_1_right_mm_read_readdatavalid,                   --                                                          .readdatavalid
			dma_comm_2_left_mm_read_address                                 => dma_comm_2_left_mm_read_address,                          --                                   dma_comm_2_left_mm_read.address
			dma_comm_2_left_mm_read_waitrequest                             => dma_comm_2_left_mm_read_waitrequest,                      --                                                          .waitrequest
			dma_comm_2_left_mm_read_byteenable                              => dma_comm_2_left_mm_read_byteenable,                       --                                                          .byteenable
			dma_comm_2_left_mm_read_read                                    => dma_comm_2_left_mm_read_read,                             --                                                          .read
			dma_comm_2_left_mm_read_readdata                                => dma_comm_2_left_mm_read_readdata,                         --                                                          .readdata
			dma_comm_2_left_mm_read_readdatavalid                           => dma_comm_2_left_mm_read_readdatavalid,                    --                                                          .readdatavalid
			dma_comm_2_right_mm_read_address                                => dma_comm_2_right_mm_read_address,                         --                                  dma_comm_2_right_mm_read.address
			dma_comm_2_right_mm_read_waitrequest                            => dma_comm_2_right_mm_read_waitrequest,                     --                                                          .waitrequest
			dma_comm_2_right_mm_read_byteenable                             => dma_comm_2_right_mm_read_byteenable,                      --                                                          .byteenable
			dma_comm_2_right_mm_read_read                                   => dma_comm_2_right_mm_read_read,                            --                                                          .read
			dma_comm_2_right_mm_read_readdata                               => dma_comm_2_right_mm_read_readdata,                        --                                                          .readdata
			dma_comm_2_right_mm_read_readdatavalid                          => dma_comm_2_right_mm_read_readdatavalid,                   --                                                          .readdatavalid
			dma_comm_3_left_mm_read_address                                 => dma_comm_3_left_mm_read_address,                          --                                   dma_comm_3_left_mm_read.address
			dma_comm_3_left_mm_read_waitrequest                             => dma_comm_3_left_mm_read_waitrequest,                      --                                                          .waitrequest
			dma_comm_3_left_mm_read_byteenable                              => dma_comm_3_left_mm_read_byteenable,                       --                                                          .byteenable
			dma_comm_3_left_mm_read_read                                    => dma_comm_3_left_mm_read_read,                             --                                                          .read
			dma_comm_3_left_mm_read_readdata                                => dma_comm_3_left_mm_read_readdata,                         --                                                          .readdata
			dma_comm_3_left_mm_read_readdatavalid                           => dma_comm_3_left_mm_read_readdatavalid,                    --                                                          .readdatavalid
			dma_comm_3_right_mm_read_address                                => dma_comm_3_right_mm_read_address,                         --                                  dma_comm_3_right_mm_read.address
			dma_comm_3_right_mm_read_waitrequest                            => dma_comm_3_right_mm_read_waitrequest,                     --                                                          .waitrequest
			dma_comm_3_right_mm_read_byteenable                             => dma_comm_3_right_mm_read_byteenable,                      --                                                          .byteenable
			dma_comm_3_right_mm_read_read                                   => dma_comm_3_right_mm_read_read,                            --                                                          .read
			dma_comm_3_right_mm_read_readdata                               => dma_comm_3_right_mm_read_readdata,                        --                                                          .readdata
			dma_comm_3_right_mm_read_readdatavalid                          => dma_comm_3_right_mm_read_readdatavalid,                   --                                                          .readdatavalid
			dma_comm_4_left_mm_read_address                                 => dma_comm_4_left_mm_read_address,                          --                                   dma_comm_4_left_mm_read.address
			dma_comm_4_left_mm_read_waitrequest                             => dma_comm_4_left_mm_read_waitrequest,                      --                                                          .waitrequest
			dma_comm_4_left_mm_read_byteenable                              => dma_comm_4_left_mm_read_byteenable,                       --                                                          .byteenable
			dma_comm_4_left_mm_read_read                                    => dma_comm_4_left_mm_read_read,                             --                                                          .read
			dma_comm_4_left_mm_read_readdata                                => dma_comm_4_left_mm_read_readdata,                         --                                                          .readdata
			dma_comm_4_left_mm_read_readdatavalid                           => dma_comm_4_left_mm_read_readdatavalid,                    --                                                          .readdatavalid
			dma_comm_4_right_mm_read_address                                => dma_comm_4_right_mm_read_address,                         --                                  dma_comm_4_right_mm_read.address
			dma_comm_4_right_mm_read_waitrequest                            => dma_comm_4_right_mm_read_waitrequest,                     --                                                          .waitrequest
			dma_comm_4_right_mm_read_byteenable                             => dma_comm_4_right_mm_read_byteenable,                      --                                                          .byteenable
			dma_comm_4_right_mm_read_read                                   => dma_comm_4_right_mm_read_read,                            --                                                          .read
			dma_comm_4_right_mm_read_readdata                               => dma_comm_4_right_mm_read_readdata,                        --                                                          .readdata
			dma_comm_4_right_mm_read_readdatavalid                          => dma_comm_4_right_mm_read_readdatavalid,                   --                                                          .readdatavalid
			dma_comm_5_left_mm_read_address                                 => dma_comm_5_left_mm_read_address,                          --                                   dma_comm_5_left_mm_read.address
			dma_comm_5_left_mm_read_waitrequest                             => dma_comm_5_left_mm_read_waitrequest,                      --                                                          .waitrequest
			dma_comm_5_left_mm_read_byteenable                              => dma_comm_5_left_mm_read_byteenable,                       --                                                          .byteenable
			dma_comm_5_left_mm_read_read                                    => dma_comm_5_left_mm_read_read,                             --                                                          .read
			dma_comm_5_left_mm_read_readdata                                => dma_comm_5_left_mm_read_readdata,                         --                                                          .readdata
			dma_comm_5_left_mm_read_readdatavalid                           => dma_comm_5_left_mm_read_readdatavalid,                    --                                                          .readdatavalid
			dma_comm_5_right_mm_read_address                                => dma_comm_5_right_mm_read_address,                         --                                  dma_comm_5_right_mm_read.address
			dma_comm_5_right_mm_read_waitrequest                            => dma_comm_5_right_mm_read_waitrequest,                     --                                                          .waitrequest
			dma_comm_5_right_mm_read_byteenable                             => dma_comm_5_right_mm_read_byteenable,                      --                                                          .byteenable
			dma_comm_5_right_mm_read_read                                   => dma_comm_5_right_mm_read_read,                            --                                                          .read
			dma_comm_5_right_mm_read_readdata                               => dma_comm_5_right_mm_read_readdata,                        --                                                          .readdata
			dma_comm_5_right_mm_read_readdatavalid                          => dma_comm_5_right_mm_read_readdatavalid,                   --                                                          .readdatavalid
			dma_comm_6_left_mm_read_address                                 => dma_comm_6_left_mm_read_address,                          --                                   dma_comm_6_left_mm_read.address
			dma_comm_6_left_mm_read_waitrequest                             => dma_comm_6_left_mm_read_waitrequest,                      --                                                          .waitrequest
			dma_comm_6_left_mm_read_byteenable                              => dma_comm_6_left_mm_read_byteenable,                       --                                                          .byteenable
			dma_comm_6_left_mm_read_read                                    => dma_comm_6_left_mm_read_read,                             --                                                          .read
			dma_comm_6_left_mm_read_readdata                                => dma_comm_6_left_mm_read_readdata,                         --                                                          .readdata
			dma_comm_6_left_mm_read_readdatavalid                           => dma_comm_6_left_mm_read_readdatavalid,                    --                                                          .readdatavalid
			dma_comm_6_right_mm_read_address                                => dma_comm_6_right_mm_read_address,                         --                                  dma_comm_6_right_mm_read.address
			dma_comm_6_right_mm_read_waitrequest                            => dma_comm_6_right_mm_read_waitrequest,                     --                                                          .waitrequest
			dma_comm_6_right_mm_read_byteenable                             => dma_comm_6_right_mm_read_byteenable,                      --                                                          .byteenable
			dma_comm_6_right_mm_read_read                                   => dma_comm_6_right_mm_read_read,                            --                                                          .read
			dma_comm_6_right_mm_read_readdata                               => dma_comm_6_right_mm_read_readdata,                        --                                                          .readdata
			dma_comm_6_right_mm_read_readdatavalid                          => dma_comm_6_right_mm_read_readdatavalid,                   --                                                          .readdatavalid
			dma_ftdi_usb3_mm_write_address                                  => dma_ftdi_usb3_mm_write_address,                           --                                    dma_ftdi_usb3_mm_write.address
			dma_ftdi_usb3_mm_write_waitrequest                              => dma_ftdi_usb3_mm_write_waitrequest,                       --                                                          .waitrequest
			dma_ftdi_usb3_mm_write_byteenable                               => dma_ftdi_usb3_mm_write_byteenable,                        --                                                          .byteenable
			dma_ftdi_usb3_mm_write_write                                    => dma_ftdi_usb3_mm_write_write,                             --                                                          .write
			dma_ftdi_usb3_mm_write_writedata                                => dma_ftdi_usb3_mm_write_writedata,                         --                                                          .writedata
			rmap_mem_nfee_comm_1_avalon_mm_rmap_master_address              => rmap_mem_nfee_comm_1_avalon_mm_rmap_master_address,       --                rmap_mem_nfee_comm_1_avalon_mm_rmap_master.address
			rmap_mem_nfee_comm_1_avalon_mm_rmap_master_waitrequest          => rmap_mem_nfee_comm_1_avalon_mm_rmap_master_waitrequest,   --                                                          .waitrequest
			rmap_mem_nfee_comm_1_avalon_mm_rmap_master_read                 => rmap_mem_nfee_comm_1_avalon_mm_rmap_master_read,          --                                                          .read
			rmap_mem_nfee_comm_1_avalon_mm_rmap_master_readdata             => rmap_mem_nfee_comm_1_avalon_mm_rmap_master_readdata,      --                                                          .readdata
			rmap_mem_nfee_comm_1_avalon_mm_rmap_master_write                => rmap_mem_nfee_comm_1_avalon_mm_rmap_master_write,         --                                                          .write
			rmap_mem_nfee_comm_1_avalon_mm_rmap_master_writedata            => rmap_mem_nfee_comm_1_avalon_mm_rmap_master_writedata,     --                                                          .writedata
			rmap_mem_nfee_comm_2_avalon_mm_rmap_master_address              => rmap_mem_nfee_comm_2_avalon_mm_rmap_master_address,       --                rmap_mem_nfee_comm_2_avalon_mm_rmap_master.address
			rmap_mem_nfee_comm_2_avalon_mm_rmap_master_waitrequest          => rmap_mem_nfee_comm_2_avalon_mm_rmap_master_waitrequest,   --                                                          .waitrequest
			rmap_mem_nfee_comm_2_avalon_mm_rmap_master_read                 => rmap_mem_nfee_comm_2_avalon_mm_rmap_master_read,          --                                                          .read
			rmap_mem_nfee_comm_2_avalon_mm_rmap_master_readdata             => rmap_mem_nfee_comm_2_avalon_mm_rmap_master_readdata,      --                                                          .readdata
			rmap_mem_nfee_comm_2_avalon_mm_rmap_master_write                => rmap_mem_nfee_comm_2_avalon_mm_rmap_master_write,         --                                                          .write
			rmap_mem_nfee_comm_2_avalon_mm_rmap_master_writedata            => rmap_mem_nfee_comm_2_avalon_mm_rmap_master_writedata,     --                                                          .writedata
			rmap_mem_nfee_comm_3_avalon_mm_rmap_master_address              => rmap_mem_nfee_comm_3_avalon_mm_rmap_master_address,       --                rmap_mem_nfee_comm_3_avalon_mm_rmap_master.address
			rmap_mem_nfee_comm_3_avalon_mm_rmap_master_waitrequest          => rmap_mem_nfee_comm_3_avalon_mm_rmap_master_waitrequest,   --                                                          .waitrequest
			rmap_mem_nfee_comm_3_avalon_mm_rmap_master_read                 => rmap_mem_nfee_comm_3_avalon_mm_rmap_master_read,          --                                                          .read
			rmap_mem_nfee_comm_3_avalon_mm_rmap_master_readdata             => rmap_mem_nfee_comm_3_avalon_mm_rmap_master_readdata,      --                                                          .readdata
			rmap_mem_nfee_comm_3_avalon_mm_rmap_master_write                => rmap_mem_nfee_comm_3_avalon_mm_rmap_master_write,         --                                                          .write
			rmap_mem_nfee_comm_3_avalon_mm_rmap_master_writedata            => rmap_mem_nfee_comm_3_avalon_mm_rmap_master_writedata,     --                                                          .writedata
			rmap_mem_nfee_comm_4_avalon_mm_rmap_master_address              => rmap_mem_nfee_comm_4_avalon_mm_rmap_master_address,       --                rmap_mem_nfee_comm_4_avalon_mm_rmap_master.address
			rmap_mem_nfee_comm_4_avalon_mm_rmap_master_waitrequest          => rmap_mem_nfee_comm_4_avalon_mm_rmap_master_waitrequest,   --                                                          .waitrequest
			rmap_mem_nfee_comm_4_avalon_mm_rmap_master_read                 => rmap_mem_nfee_comm_4_avalon_mm_rmap_master_read,          --                                                          .read
			rmap_mem_nfee_comm_4_avalon_mm_rmap_master_readdata             => rmap_mem_nfee_comm_4_avalon_mm_rmap_master_readdata,      --                                                          .readdata
			rmap_mem_nfee_comm_4_avalon_mm_rmap_master_write                => rmap_mem_nfee_comm_4_avalon_mm_rmap_master_write,         --                                                          .write
			rmap_mem_nfee_comm_4_avalon_mm_rmap_master_writedata            => rmap_mem_nfee_comm_4_avalon_mm_rmap_master_writedata,     --                                                          .writedata
			rmap_mem_nfee_comm_5_avalon_mm_rmap_master_address              => rmap_mem_nfee_comm_5_avalon_mm_rmap_master_address,       --                rmap_mem_nfee_comm_5_avalon_mm_rmap_master.address
			rmap_mem_nfee_comm_5_avalon_mm_rmap_master_waitrequest          => rmap_mem_nfee_comm_5_avalon_mm_rmap_master_waitrequest,   --                                                          .waitrequest
			rmap_mem_nfee_comm_5_avalon_mm_rmap_master_read                 => rmap_mem_nfee_comm_5_avalon_mm_rmap_master_read,          --                                                          .read
			rmap_mem_nfee_comm_5_avalon_mm_rmap_master_readdata             => rmap_mem_nfee_comm_5_avalon_mm_rmap_master_readdata,      --                                                          .readdata
			rmap_mem_nfee_comm_5_avalon_mm_rmap_master_write                => rmap_mem_nfee_comm_5_avalon_mm_rmap_master_write,         --                                                          .write
			rmap_mem_nfee_comm_5_avalon_mm_rmap_master_writedata            => rmap_mem_nfee_comm_5_avalon_mm_rmap_master_writedata,     --                                                          .writedata
			rmap_mem_nfee_comm_6_avalon_mm_rmap_master_address              => rmap_mem_nfee_comm_6_avalon_mm_rmap_master_address,       --                rmap_mem_nfee_comm_6_avalon_mm_rmap_master.address
			rmap_mem_nfee_comm_6_avalon_mm_rmap_master_waitrequest          => rmap_mem_nfee_comm_6_avalon_mm_rmap_master_waitrequest,   --                                                          .waitrequest
			rmap_mem_nfee_comm_6_avalon_mm_rmap_master_read                 => rmap_mem_nfee_comm_6_avalon_mm_rmap_master_read,          --                                                          .read
			rmap_mem_nfee_comm_6_avalon_mm_rmap_master_readdata             => rmap_mem_nfee_comm_6_avalon_mm_rmap_master_readdata,      --                                                          .readdata
			rmap_mem_nfee_comm_6_avalon_mm_rmap_master_write                => rmap_mem_nfee_comm_6_avalon_mm_rmap_master_write,         --                                                          .write
			rmap_mem_nfee_comm_6_avalon_mm_rmap_master_writedata            => rmap_mem_nfee_comm_6_avalon_mm_rmap_master_writedata,     --                                                          .writedata
			m1_clock_bridge_s0_address                                      => mm_interconnect_0_m1_clock_bridge_s0_address,             --                                        m1_clock_bridge_s0.address
			m1_clock_bridge_s0_write                                        => mm_interconnect_0_m1_clock_bridge_s0_write,               --                                                          .write
			m1_clock_bridge_s0_read                                         => mm_interconnect_0_m1_clock_bridge_s0_read,                --                                                          .read
			m1_clock_bridge_s0_readdata                                     => mm_interconnect_0_m1_clock_bridge_s0_readdata,            --                                                          .readdata
			m1_clock_bridge_s0_writedata                                    => mm_interconnect_0_m1_clock_bridge_s0_writedata,           --                                                          .writedata
			m1_clock_bridge_s0_burstcount                                   => mm_interconnect_0_m1_clock_bridge_s0_burstcount,          --                                                          .burstcount
			m1_clock_bridge_s0_byteenable                                   => mm_interconnect_0_m1_clock_bridge_s0_byteenable,          --                                                          .byteenable
			m1_clock_bridge_s0_readdatavalid                                => mm_interconnect_0_m1_clock_bridge_s0_readdatavalid,       --                                                          .readdatavalid
			m1_clock_bridge_s0_waitrequest                                  => mm_interconnect_0_m1_clock_bridge_s0_waitrequest,         --                                                          .waitrequest
			m1_clock_bridge_s0_debugaccess                                  => mm_interconnect_0_m1_clock_bridge_s0_debugaccess,         --                                                          .debugaccess
			m2_ddr2_memory_avl_address                                      => mm_interconnect_0_m2_ddr2_memory_avl_address,             --                                        m2_ddr2_memory_avl.address
			m2_ddr2_memory_avl_write                                        => mm_interconnect_0_m2_ddr2_memory_avl_write,               --                                                          .write
			m2_ddr2_memory_avl_read                                         => mm_interconnect_0_m2_ddr2_memory_avl_read,                --                                                          .read
			m2_ddr2_memory_avl_readdata                                     => mm_interconnect_0_m2_ddr2_memory_avl_readdata,            --                                                          .readdata
			m2_ddr2_memory_avl_writedata                                    => mm_interconnect_0_m2_ddr2_memory_avl_writedata,           --                                                          .writedata
			m2_ddr2_memory_avl_beginbursttransfer                           => mm_interconnect_0_m2_ddr2_memory_avl_beginbursttransfer,  --                                                          .beginbursttransfer
			m2_ddr2_memory_avl_burstcount                                   => mm_interconnect_0_m2_ddr2_memory_avl_burstcount,          --                                                          .burstcount
			m2_ddr2_memory_avl_byteenable                                   => mm_interconnect_0_m2_ddr2_memory_avl_byteenable,          --                                                          .byteenable
			m2_ddr2_memory_avl_readdatavalid                                => mm_interconnect_0_m2_ddr2_memory_avl_readdatavalid,       --                                                          .readdatavalid
			m2_ddr2_memory_avl_waitrequest                                  => mm_interconnect_0_m2_ddr2_memory_avl_inv                  --                                                          .waitrequest
		);

	mm_interconnect_1 : component MebX_Qsys_Project_mm_interconnect_1
		port map (
			clk_100_clk_clk                                             => m2_ddr2_memory_afi_half_clk_clk,                                            --                                           clk_100_clk.clk
			ext_flash_reset_reset_bridge_in_reset_reset                 => rst_controller_010_reset_out_reset,                                         --                 ext_flash_reset_reset_bridge_in_reset.reset
			jtag_uart_0_reset_reset_bridge_in_reset_reset               => rst_controller_008_reset_out_reset,                                         --               jtag_uart_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset              => rst_controller_012_reset_out_reset,                                         --              nios2_gen2_0_reset_reset_bridge_in_reset.reset
			rmap_mem_nfee_comm_1_reset_sink_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                                         -- rmap_mem_nfee_comm_1_reset_sink_reset_bridge_in_reset.reset
			rmap_mem_nfee_comm_2_reset_sink_reset_bridge_in_reset_reset => rst_controller_003_reset_out_reset,                                         -- rmap_mem_nfee_comm_2_reset_sink_reset_bridge_in_reset.reset
			rmap_mem_nfee_comm_3_reset_sink_reset_bridge_in_reset_reset => rst_controller_004_reset_out_reset,                                         -- rmap_mem_nfee_comm_3_reset_sink_reset_bridge_in_reset.reset
			rmap_mem_nfee_comm_4_reset_sink_reset_bridge_in_reset_reset => rst_controller_005_reset_out_reset,                                         -- rmap_mem_nfee_comm_4_reset_sink_reset_bridge_in_reset.reset
			rmap_mem_nfee_comm_5_reset_sink_reset_bridge_in_reset_reset => rst_controller_006_reset_out_reset,                                         -- rmap_mem_nfee_comm_5_reset_sink_reset_bridge_in_reset.reset
			rmap_mem_nfee_comm_6_reset_sink_reset_bridge_in_reset_reset => rst_controller_007_reset_out_reset,                                         -- rmap_mem_nfee_comm_6_reset_sink_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                            => nios2_gen2_0_data_master_address,                                           --                              nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                        => nios2_gen2_0_data_master_waitrequest,                                       --                                                      .waitrequest
			nios2_gen2_0_data_master_byteenable                         => nios2_gen2_0_data_master_byteenable,                                        --                                                      .byteenable
			nios2_gen2_0_data_master_read                               => nios2_gen2_0_data_master_read,                                              --                                                      .read
			nios2_gen2_0_data_master_readdata                           => nios2_gen2_0_data_master_readdata,                                          --                                                      .readdata
			nios2_gen2_0_data_master_write                              => nios2_gen2_0_data_master_write,                                             --                                                      .write
			nios2_gen2_0_data_master_writedata                          => nios2_gen2_0_data_master_writedata,                                         --                                                      .writedata
			nios2_gen2_0_data_master_debugaccess                        => nios2_gen2_0_data_master_debugaccess,                                       --                                                      .debugaccess
			nios2_gen2_0_instruction_master_address                     => nios2_gen2_0_instruction_master_address,                                    --                       nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest                 => nios2_gen2_0_instruction_master_waitrequest,                                --                                                      .waitrequest
			nios2_gen2_0_instruction_master_burstcount                  => nios2_gen2_0_instruction_master_burstcount,                                 --                                                      .burstcount
			nios2_gen2_0_instruction_master_read                        => nios2_gen2_0_instruction_master_read,                                       --                                                      .read
			nios2_gen2_0_instruction_master_readdata                    => nios2_gen2_0_instruction_master_readdata,                                   --                                                      .readdata
			nios2_gen2_0_instruction_master_readdatavalid               => nios2_gen2_0_instruction_master_readdatavalid,                              --                                                      .readdatavalid
			clock_bridge_afi_50_s0_address                              => mm_interconnect_1_clock_bridge_afi_50_s0_address,                           --                                clock_bridge_afi_50_s0.address
			clock_bridge_afi_50_s0_write                                => mm_interconnect_1_clock_bridge_afi_50_s0_write,                             --                                                      .write
			clock_bridge_afi_50_s0_read                                 => mm_interconnect_1_clock_bridge_afi_50_s0_read,                              --                                                      .read
			clock_bridge_afi_50_s0_readdata                             => mm_interconnect_1_clock_bridge_afi_50_s0_readdata,                          --                                                      .readdata
			clock_bridge_afi_50_s0_writedata                            => mm_interconnect_1_clock_bridge_afi_50_s0_writedata,                         --                                                      .writedata
			clock_bridge_afi_50_s0_burstcount                           => mm_interconnect_1_clock_bridge_afi_50_s0_burstcount,                        --                                                      .burstcount
			clock_bridge_afi_50_s0_byteenable                           => mm_interconnect_1_clock_bridge_afi_50_s0_byteenable,                        --                                                      .byteenable
			clock_bridge_afi_50_s0_readdatavalid                        => mm_interconnect_1_clock_bridge_afi_50_s0_readdatavalid,                     --                                                      .readdatavalid
			clock_bridge_afi_50_s0_waitrequest                          => mm_interconnect_1_clock_bridge_afi_50_s0_waitrequest,                       --                                                      .waitrequest
			clock_bridge_afi_50_s0_debugaccess                          => mm_interconnect_1_clock_bridge_afi_50_s0_debugaccess,                       --                                                      .debugaccess
			COMM_Pedreiro_v1_01_A_avalon_slave_windowing_address        => mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_address,     --          COMM_Pedreiro_v1_01_A_avalon_slave_windowing.address
			COMM_Pedreiro_v1_01_A_avalon_slave_windowing_write          => mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_write,       --                                                      .write
			COMM_Pedreiro_v1_01_A_avalon_slave_windowing_read           => mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_read,        --                                                      .read
			COMM_Pedreiro_v1_01_A_avalon_slave_windowing_readdata       => mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_readdata,    --                                                      .readdata
			COMM_Pedreiro_v1_01_A_avalon_slave_windowing_writedata      => mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_writedata,   --                                                      .writedata
			COMM_Pedreiro_v1_01_A_avalon_slave_windowing_byteenable     => mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_byteenable,  --                                                      .byteenable
			COMM_Pedreiro_v1_01_A_avalon_slave_windowing_waitrequest    => mm_interconnect_1_comm_pedreiro_v1_01_a_avalon_slave_windowing_waitrequest, --                                                      .waitrequest
			COMM_Pedreiro_v1_01_B_avalon_slave_windowing_address        => mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_address,     --          COMM_Pedreiro_v1_01_B_avalon_slave_windowing.address
			COMM_Pedreiro_v1_01_B_avalon_slave_windowing_write          => mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_write,       --                                                      .write
			COMM_Pedreiro_v1_01_B_avalon_slave_windowing_read           => mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_read,        --                                                      .read
			COMM_Pedreiro_v1_01_B_avalon_slave_windowing_readdata       => mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_readdata,    --                                                      .readdata
			COMM_Pedreiro_v1_01_B_avalon_slave_windowing_writedata      => mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_writedata,   --                                                      .writedata
			COMM_Pedreiro_v1_01_B_avalon_slave_windowing_byteenable     => mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_byteenable,  --                                                      .byteenable
			COMM_Pedreiro_v1_01_B_avalon_slave_windowing_waitrequest    => mm_interconnect_1_comm_pedreiro_v1_01_b_avalon_slave_windowing_waitrequest, --                                                      .waitrequest
			COMM_Pedreiro_v1_01_C_avalon_slave_windowing_address        => mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_address,     --          COMM_Pedreiro_v1_01_C_avalon_slave_windowing.address
			COMM_Pedreiro_v1_01_C_avalon_slave_windowing_write          => mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_write,       --                                                      .write
			COMM_Pedreiro_v1_01_C_avalon_slave_windowing_read           => mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_read,        --                                                      .read
			COMM_Pedreiro_v1_01_C_avalon_slave_windowing_readdata       => mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_readdata,    --                                                      .readdata
			COMM_Pedreiro_v1_01_C_avalon_slave_windowing_writedata      => mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_writedata,   --                                                      .writedata
			COMM_Pedreiro_v1_01_C_avalon_slave_windowing_byteenable     => mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_byteenable,  --                                                      .byteenable
			COMM_Pedreiro_v1_01_C_avalon_slave_windowing_waitrequest    => mm_interconnect_1_comm_pedreiro_v1_01_c_avalon_slave_windowing_waitrequest, --                                                      .waitrequest
			COMM_Pedreiro_v1_01_D_avalon_slave_windowing_address        => mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_address,     --          COMM_Pedreiro_v1_01_D_avalon_slave_windowing.address
			COMM_Pedreiro_v1_01_D_avalon_slave_windowing_write          => mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_write,       --                                                      .write
			COMM_Pedreiro_v1_01_D_avalon_slave_windowing_read           => mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_read,        --                                                      .read
			COMM_Pedreiro_v1_01_D_avalon_slave_windowing_readdata       => mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_readdata,    --                                                      .readdata
			COMM_Pedreiro_v1_01_D_avalon_slave_windowing_writedata      => mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_writedata,   --                                                      .writedata
			COMM_Pedreiro_v1_01_D_avalon_slave_windowing_byteenable     => mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_byteenable,  --                                                      .byteenable
			COMM_Pedreiro_v1_01_D_avalon_slave_windowing_waitrequest    => mm_interconnect_1_comm_pedreiro_v1_01_d_avalon_slave_windowing_waitrequest, --                                                      .waitrequest
			COMM_Pedreiro_v1_01_E_avalon_slave_windowing_address        => mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_address,     --          COMM_Pedreiro_v1_01_E_avalon_slave_windowing.address
			COMM_Pedreiro_v1_01_E_avalon_slave_windowing_write          => mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_write,       --                                                      .write
			COMM_Pedreiro_v1_01_E_avalon_slave_windowing_read           => mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_read,        --                                                      .read
			COMM_Pedreiro_v1_01_E_avalon_slave_windowing_readdata       => mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_readdata,    --                                                      .readdata
			COMM_Pedreiro_v1_01_E_avalon_slave_windowing_writedata      => mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_writedata,   --                                                      .writedata
			COMM_Pedreiro_v1_01_E_avalon_slave_windowing_byteenable     => mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_byteenable,  --                                                      .byteenable
			COMM_Pedreiro_v1_01_E_avalon_slave_windowing_waitrequest    => mm_interconnect_1_comm_pedreiro_v1_01_e_avalon_slave_windowing_waitrequest, --                                                      .waitrequest
			COMM_Pedreiro_v1_01_F_avalon_slave_windowing_address        => mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_address,     --          COMM_Pedreiro_v1_01_F_avalon_slave_windowing.address
			COMM_Pedreiro_v1_01_F_avalon_slave_windowing_write          => mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_write,       --                                                      .write
			COMM_Pedreiro_v1_01_F_avalon_slave_windowing_read           => mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_read,        --                                                      .read
			COMM_Pedreiro_v1_01_F_avalon_slave_windowing_readdata       => mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_readdata,    --                                                      .readdata
			COMM_Pedreiro_v1_01_F_avalon_slave_windowing_writedata      => mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_writedata,   --                                                      .writedata
			COMM_Pedreiro_v1_01_F_avalon_slave_windowing_byteenable     => mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_byteenable,  --                                                      .byteenable
			COMM_Pedreiro_v1_01_F_avalon_slave_windowing_waitrequest    => mm_interconnect_1_comm_pedreiro_v1_01_f_avalon_slave_windowing_waitrequest, --                                                      .waitrequest
			ddr2_address_span_extender_cntl_write                       => mm_interconnect_1_ddr2_address_span_extender_cntl_write,                    --                       ddr2_address_span_extender_cntl.write
			ddr2_address_span_extender_cntl_read                        => mm_interconnect_1_ddr2_address_span_extender_cntl_read,                     --                                                      .read
			ddr2_address_span_extender_cntl_readdata                    => mm_interconnect_1_ddr2_address_span_extender_cntl_readdata,                 --                                                      .readdata
			ddr2_address_span_extender_cntl_writedata                   => mm_interconnect_1_ddr2_address_span_extender_cntl_writedata,                --                                                      .writedata
			ddr2_address_span_extender_cntl_byteenable                  => mm_interconnect_1_ddr2_address_span_extender_cntl_byteenable,               --                                                      .byteenable
			ddr2_address_span_extender_windowed_slave_address           => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_address,        --             ddr2_address_span_extender_windowed_slave.address
			ddr2_address_span_extender_windowed_slave_write             => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_write,          --                                                      .write
			ddr2_address_span_extender_windowed_slave_read              => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_read,           --                                                      .read
			ddr2_address_span_extender_windowed_slave_readdata          => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdata,       --                                                      .readdata
			ddr2_address_span_extender_windowed_slave_writedata         => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_writedata,      --                                                      .writedata
			ddr2_address_span_extender_windowed_slave_burstcount        => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_burstcount,     --                                                      .burstcount
			ddr2_address_span_extender_windowed_slave_byteenable        => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_byteenable,     --                                                      .byteenable
			ddr2_address_span_extender_windowed_slave_readdatavalid     => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_readdatavalid,  --                                                      .readdatavalid
			ddr2_address_span_extender_windowed_slave_waitrequest       => mm_interconnect_1_ddr2_address_span_extender_windowed_slave_waitrequest,    --                                                      .waitrequest
			dma_comm_1_left_csr_address                                 => mm_interconnect_1_dma_comm_1_left_csr_address,                              --                                   dma_comm_1_left_csr.address
			dma_comm_1_left_csr_write                                   => mm_interconnect_1_dma_comm_1_left_csr_write,                                --                                                      .write
			dma_comm_1_left_csr_read                                    => mm_interconnect_1_dma_comm_1_left_csr_read,                                 --                                                      .read
			dma_comm_1_left_csr_readdata                                => mm_interconnect_1_dma_comm_1_left_csr_readdata,                             --                                                      .readdata
			dma_comm_1_left_csr_writedata                               => mm_interconnect_1_dma_comm_1_left_csr_writedata,                            --                                                      .writedata
			dma_comm_1_left_csr_byteenable                              => mm_interconnect_1_dma_comm_1_left_csr_byteenable,                           --                                                      .byteenable
			dma_comm_1_left_descriptor_slave_write                      => mm_interconnect_1_dma_comm_1_left_descriptor_slave_write,                   --                      dma_comm_1_left_descriptor_slave.write
			dma_comm_1_left_descriptor_slave_writedata                  => mm_interconnect_1_dma_comm_1_left_descriptor_slave_writedata,               --                                                      .writedata
			dma_comm_1_left_descriptor_slave_byteenable                 => mm_interconnect_1_dma_comm_1_left_descriptor_slave_byteenable,              --                                                      .byteenable
			dma_comm_1_left_descriptor_slave_waitrequest                => mm_interconnect_1_dma_comm_1_left_descriptor_slave_waitrequest,             --                                                      .waitrequest
			dma_comm_1_right_csr_address                                => mm_interconnect_1_dma_comm_1_right_csr_address,                             --                                  dma_comm_1_right_csr.address
			dma_comm_1_right_csr_write                                  => mm_interconnect_1_dma_comm_1_right_csr_write,                               --                                                      .write
			dma_comm_1_right_csr_read                                   => mm_interconnect_1_dma_comm_1_right_csr_read,                                --                                                      .read
			dma_comm_1_right_csr_readdata                               => mm_interconnect_1_dma_comm_1_right_csr_readdata,                            --                                                      .readdata
			dma_comm_1_right_csr_writedata                              => mm_interconnect_1_dma_comm_1_right_csr_writedata,                           --                                                      .writedata
			dma_comm_1_right_csr_byteenable                             => mm_interconnect_1_dma_comm_1_right_csr_byteenable,                          --                                                      .byteenable
			dma_comm_1_right_descriptor_slave_write                     => mm_interconnect_1_dma_comm_1_right_descriptor_slave_write,                  --                     dma_comm_1_right_descriptor_slave.write
			dma_comm_1_right_descriptor_slave_writedata                 => mm_interconnect_1_dma_comm_1_right_descriptor_slave_writedata,              --                                                      .writedata
			dma_comm_1_right_descriptor_slave_byteenable                => mm_interconnect_1_dma_comm_1_right_descriptor_slave_byteenable,             --                                                      .byteenable
			dma_comm_1_right_descriptor_slave_waitrequest               => mm_interconnect_1_dma_comm_1_right_descriptor_slave_waitrequest,            --                                                      .waitrequest
			dma_comm_2_left_csr_address                                 => mm_interconnect_1_dma_comm_2_left_csr_address,                              --                                   dma_comm_2_left_csr.address
			dma_comm_2_left_csr_write                                   => mm_interconnect_1_dma_comm_2_left_csr_write,                                --                                                      .write
			dma_comm_2_left_csr_read                                    => mm_interconnect_1_dma_comm_2_left_csr_read,                                 --                                                      .read
			dma_comm_2_left_csr_readdata                                => mm_interconnect_1_dma_comm_2_left_csr_readdata,                             --                                                      .readdata
			dma_comm_2_left_csr_writedata                               => mm_interconnect_1_dma_comm_2_left_csr_writedata,                            --                                                      .writedata
			dma_comm_2_left_csr_byteenable                              => mm_interconnect_1_dma_comm_2_left_csr_byteenable,                           --                                                      .byteenable
			dma_comm_2_left_descriptor_slave_write                      => mm_interconnect_1_dma_comm_2_left_descriptor_slave_write,                   --                      dma_comm_2_left_descriptor_slave.write
			dma_comm_2_left_descriptor_slave_writedata                  => mm_interconnect_1_dma_comm_2_left_descriptor_slave_writedata,               --                                                      .writedata
			dma_comm_2_left_descriptor_slave_byteenable                 => mm_interconnect_1_dma_comm_2_left_descriptor_slave_byteenable,              --                                                      .byteenable
			dma_comm_2_left_descriptor_slave_waitrequest                => mm_interconnect_1_dma_comm_2_left_descriptor_slave_waitrequest,             --                                                      .waitrequest
			dma_comm_2_right_csr_address                                => mm_interconnect_1_dma_comm_2_right_csr_address,                             --                                  dma_comm_2_right_csr.address
			dma_comm_2_right_csr_write                                  => mm_interconnect_1_dma_comm_2_right_csr_write,                               --                                                      .write
			dma_comm_2_right_csr_read                                   => mm_interconnect_1_dma_comm_2_right_csr_read,                                --                                                      .read
			dma_comm_2_right_csr_readdata                               => mm_interconnect_1_dma_comm_2_right_csr_readdata,                            --                                                      .readdata
			dma_comm_2_right_csr_writedata                              => mm_interconnect_1_dma_comm_2_right_csr_writedata,                           --                                                      .writedata
			dma_comm_2_right_csr_byteenable                             => mm_interconnect_1_dma_comm_2_right_csr_byteenable,                          --                                                      .byteenable
			dma_comm_2_right_descriptor_slave_write                     => mm_interconnect_1_dma_comm_2_right_descriptor_slave_write,                  --                     dma_comm_2_right_descriptor_slave.write
			dma_comm_2_right_descriptor_slave_writedata                 => mm_interconnect_1_dma_comm_2_right_descriptor_slave_writedata,              --                                                      .writedata
			dma_comm_2_right_descriptor_slave_byteenable                => mm_interconnect_1_dma_comm_2_right_descriptor_slave_byteenable,             --                                                      .byteenable
			dma_comm_2_right_descriptor_slave_waitrequest               => mm_interconnect_1_dma_comm_2_right_descriptor_slave_waitrequest,            --                                                      .waitrequest
			dma_comm_3_left_csr_address                                 => mm_interconnect_1_dma_comm_3_left_csr_address,                              --                                   dma_comm_3_left_csr.address
			dma_comm_3_left_csr_write                                   => mm_interconnect_1_dma_comm_3_left_csr_write,                                --                                                      .write
			dma_comm_3_left_csr_read                                    => mm_interconnect_1_dma_comm_3_left_csr_read,                                 --                                                      .read
			dma_comm_3_left_csr_readdata                                => mm_interconnect_1_dma_comm_3_left_csr_readdata,                             --                                                      .readdata
			dma_comm_3_left_csr_writedata                               => mm_interconnect_1_dma_comm_3_left_csr_writedata,                            --                                                      .writedata
			dma_comm_3_left_csr_byteenable                              => mm_interconnect_1_dma_comm_3_left_csr_byteenable,                           --                                                      .byteenable
			dma_comm_3_left_descriptor_slave_write                      => mm_interconnect_1_dma_comm_3_left_descriptor_slave_write,                   --                      dma_comm_3_left_descriptor_slave.write
			dma_comm_3_left_descriptor_slave_writedata                  => mm_interconnect_1_dma_comm_3_left_descriptor_slave_writedata,               --                                                      .writedata
			dma_comm_3_left_descriptor_slave_byteenable                 => mm_interconnect_1_dma_comm_3_left_descriptor_slave_byteenable,              --                                                      .byteenable
			dma_comm_3_left_descriptor_slave_waitrequest                => mm_interconnect_1_dma_comm_3_left_descriptor_slave_waitrequest,             --                                                      .waitrequest
			dma_comm_3_right_csr_address                                => mm_interconnect_1_dma_comm_3_right_csr_address,                             --                                  dma_comm_3_right_csr.address
			dma_comm_3_right_csr_write                                  => mm_interconnect_1_dma_comm_3_right_csr_write,                               --                                                      .write
			dma_comm_3_right_csr_read                                   => mm_interconnect_1_dma_comm_3_right_csr_read,                                --                                                      .read
			dma_comm_3_right_csr_readdata                               => mm_interconnect_1_dma_comm_3_right_csr_readdata,                            --                                                      .readdata
			dma_comm_3_right_csr_writedata                              => mm_interconnect_1_dma_comm_3_right_csr_writedata,                           --                                                      .writedata
			dma_comm_3_right_csr_byteenable                             => mm_interconnect_1_dma_comm_3_right_csr_byteenable,                          --                                                      .byteenable
			dma_comm_3_right_descriptor_slave_write                     => mm_interconnect_1_dma_comm_3_right_descriptor_slave_write,                  --                     dma_comm_3_right_descriptor_slave.write
			dma_comm_3_right_descriptor_slave_writedata                 => mm_interconnect_1_dma_comm_3_right_descriptor_slave_writedata,              --                                                      .writedata
			dma_comm_3_right_descriptor_slave_byteenable                => mm_interconnect_1_dma_comm_3_right_descriptor_slave_byteenable,             --                                                      .byteenable
			dma_comm_3_right_descriptor_slave_waitrequest               => mm_interconnect_1_dma_comm_3_right_descriptor_slave_waitrequest,            --                                                      .waitrequest
			dma_comm_4_left_csr_address                                 => mm_interconnect_1_dma_comm_4_left_csr_address,                              --                                   dma_comm_4_left_csr.address
			dma_comm_4_left_csr_write                                   => mm_interconnect_1_dma_comm_4_left_csr_write,                                --                                                      .write
			dma_comm_4_left_csr_read                                    => mm_interconnect_1_dma_comm_4_left_csr_read,                                 --                                                      .read
			dma_comm_4_left_csr_readdata                                => mm_interconnect_1_dma_comm_4_left_csr_readdata,                             --                                                      .readdata
			dma_comm_4_left_csr_writedata                               => mm_interconnect_1_dma_comm_4_left_csr_writedata,                            --                                                      .writedata
			dma_comm_4_left_csr_byteenable                              => mm_interconnect_1_dma_comm_4_left_csr_byteenable,                           --                                                      .byteenable
			dma_comm_4_left_descriptor_slave_write                      => mm_interconnect_1_dma_comm_4_left_descriptor_slave_write,                   --                      dma_comm_4_left_descriptor_slave.write
			dma_comm_4_left_descriptor_slave_writedata                  => mm_interconnect_1_dma_comm_4_left_descriptor_slave_writedata,               --                                                      .writedata
			dma_comm_4_left_descriptor_slave_byteenable                 => mm_interconnect_1_dma_comm_4_left_descriptor_slave_byteenable,              --                                                      .byteenable
			dma_comm_4_left_descriptor_slave_waitrequest                => mm_interconnect_1_dma_comm_4_left_descriptor_slave_waitrequest,             --                                                      .waitrequest
			dma_comm_4_right_csr_address                                => mm_interconnect_1_dma_comm_4_right_csr_address,                             --                                  dma_comm_4_right_csr.address
			dma_comm_4_right_csr_write                                  => mm_interconnect_1_dma_comm_4_right_csr_write,                               --                                                      .write
			dma_comm_4_right_csr_read                                   => mm_interconnect_1_dma_comm_4_right_csr_read,                                --                                                      .read
			dma_comm_4_right_csr_readdata                               => mm_interconnect_1_dma_comm_4_right_csr_readdata,                            --                                                      .readdata
			dma_comm_4_right_csr_writedata                              => mm_interconnect_1_dma_comm_4_right_csr_writedata,                           --                                                      .writedata
			dma_comm_4_right_csr_byteenable                             => mm_interconnect_1_dma_comm_4_right_csr_byteenable,                          --                                                      .byteenable
			dma_comm_4_right_descriptor_slave_write                     => mm_interconnect_1_dma_comm_4_right_descriptor_slave_write,                  --                     dma_comm_4_right_descriptor_slave.write
			dma_comm_4_right_descriptor_slave_writedata                 => mm_interconnect_1_dma_comm_4_right_descriptor_slave_writedata,              --                                                      .writedata
			dma_comm_4_right_descriptor_slave_byteenable                => mm_interconnect_1_dma_comm_4_right_descriptor_slave_byteenable,             --                                                      .byteenable
			dma_comm_4_right_descriptor_slave_waitrequest               => mm_interconnect_1_dma_comm_4_right_descriptor_slave_waitrequest,            --                                                      .waitrequest
			dma_comm_5_left_csr_address                                 => mm_interconnect_1_dma_comm_5_left_csr_address,                              --                                   dma_comm_5_left_csr.address
			dma_comm_5_left_csr_write                                   => mm_interconnect_1_dma_comm_5_left_csr_write,                                --                                                      .write
			dma_comm_5_left_csr_read                                    => mm_interconnect_1_dma_comm_5_left_csr_read,                                 --                                                      .read
			dma_comm_5_left_csr_readdata                                => mm_interconnect_1_dma_comm_5_left_csr_readdata,                             --                                                      .readdata
			dma_comm_5_left_csr_writedata                               => mm_interconnect_1_dma_comm_5_left_csr_writedata,                            --                                                      .writedata
			dma_comm_5_left_csr_byteenable                              => mm_interconnect_1_dma_comm_5_left_csr_byteenable,                           --                                                      .byteenable
			dma_comm_5_left_descriptor_slave_write                      => mm_interconnect_1_dma_comm_5_left_descriptor_slave_write,                   --                      dma_comm_5_left_descriptor_slave.write
			dma_comm_5_left_descriptor_slave_writedata                  => mm_interconnect_1_dma_comm_5_left_descriptor_slave_writedata,               --                                                      .writedata
			dma_comm_5_left_descriptor_slave_byteenable                 => mm_interconnect_1_dma_comm_5_left_descriptor_slave_byteenable,              --                                                      .byteenable
			dma_comm_5_left_descriptor_slave_waitrequest                => mm_interconnect_1_dma_comm_5_left_descriptor_slave_waitrequest,             --                                                      .waitrequest
			dma_comm_5_right_csr_address                                => mm_interconnect_1_dma_comm_5_right_csr_address,                             --                                  dma_comm_5_right_csr.address
			dma_comm_5_right_csr_write                                  => mm_interconnect_1_dma_comm_5_right_csr_write,                               --                                                      .write
			dma_comm_5_right_csr_read                                   => mm_interconnect_1_dma_comm_5_right_csr_read,                                --                                                      .read
			dma_comm_5_right_csr_readdata                               => mm_interconnect_1_dma_comm_5_right_csr_readdata,                            --                                                      .readdata
			dma_comm_5_right_csr_writedata                              => mm_interconnect_1_dma_comm_5_right_csr_writedata,                           --                                                      .writedata
			dma_comm_5_right_csr_byteenable                             => mm_interconnect_1_dma_comm_5_right_csr_byteenable,                          --                                                      .byteenable
			dma_comm_5_right_descriptor_slave_write                     => mm_interconnect_1_dma_comm_5_right_descriptor_slave_write,                  --                     dma_comm_5_right_descriptor_slave.write
			dma_comm_5_right_descriptor_slave_writedata                 => mm_interconnect_1_dma_comm_5_right_descriptor_slave_writedata,              --                                                      .writedata
			dma_comm_5_right_descriptor_slave_byteenable                => mm_interconnect_1_dma_comm_5_right_descriptor_slave_byteenable,             --                                                      .byteenable
			dma_comm_5_right_descriptor_slave_waitrequest               => mm_interconnect_1_dma_comm_5_right_descriptor_slave_waitrequest,            --                                                      .waitrequest
			dma_comm_6_left_csr_address                                 => mm_interconnect_1_dma_comm_6_left_csr_address,                              --                                   dma_comm_6_left_csr.address
			dma_comm_6_left_csr_write                                   => mm_interconnect_1_dma_comm_6_left_csr_write,                                --                                                      .write
			dma_comm_6_left_csr_read                                    => mm_interconnect_1_dma_comm_6_left_csr_read,                                 --                                                      .read
			dma_comm_6_left_csr_readdata                                => mm_interconnect_1_dma_comm_6_left_csr_readdata,                             --                                                      .readdata
			dma_comm_6_left_csr_writedata                               => mm_interconnect_1_dma_comm_6_left_csr_writedata,                            --                                                      .writedata
			dma_comm_6_left_csr_byteenable                              => mm_interconnect_1_dma_comm_6_left_csr_byteenable,                           --                                                      .byteenable
			dma_comm_6_left_descriptor_slave_write                      => mm_interconnect_1_dma_comm_6_left_descriptor_slave_write,                   --                      dma_comm_6_left_descriptor_slave.write
			dma_comm_6_left_descriptor_slave_writedata                  => mm_interconnect_1_dma_comm_6_left_descriptor_slave_writedata,               --                                                      .writedata
			dma_comm_6_left_descriptor_slave_byteenable                 => mm_interconnect_1_dma_comm_6_left_descriptor_slave_byteenable,              --                                                      .byteenable
			dma_comm_6_left_descriptor_slave_waitrequest                => mm_interconnect_1_dma_comm_6_left_descriptor_slave_waitrequest,             --                                                      .waitrequest
			dma_comm_6_right_csr_address                                => mm_interconnect_1_dma_comm_6_right_csr_address,                             --                                  dma_comm_6_right_csr.address
			dma_comm_6_right_csr_write                                  => mm_interconnect_1_dma_comm_6_right_csr_write,                               --                                                      .write
			dma_comm_6_right_csr_read                                   => mm_interconnect_1_dma_comm_6_right_csr_read,                                --                                                      .read
			dma_comm_6_right_csr_readdata                               => mm_interconnect_1_dma_comm_6_right_csr_readdata,                            --                                                      .readdata
			dma_comm_6_right_csr_writedata                              => mm_interconnect_1_dma_comm_6_right_csr_writedata,                           --                                                      .writedata
			dma_comm_6_right_csr_byteenable                             => mm_interconnect_1_dma_comm_6_right_csr_byteenable,                          --                                                      .byteenable
			dma_comm_6_right_descriptor_slave_write                     => mm_interconnect_1_dma_comm_6_right_descriptor_slave_write,                  --                     dma_comm_6_right_descriptor_slave.write
			dma_comm_6_right_descriptor_slave_writedata                 => mm_interconnect_1_dma_comm_6_right_descriptor_slave_writedata,              --                                                      .writedata
			dma_comm_6_right_descriptor_slave_byteenable                => mm_interconnect_1_dma_comm_6_right_descriptor_slave_byteenable,             --                                                      .byteenable
			dma_comm_6_right_descriptor_slave_waitrequest               => mm_interconnect_1_dma_comm_6_right_descriptor_slave_waitrequest,            --                                                      .waitrequest
			dma_ftdi_usb3_csr_address                                   => mm_interconnect_1_dma_ftdi_usb3_csr_address,                                --                                     dma_ftdi_usb3_csr.address
			dma_ftdi_usb3_csr_write                                     => mm_interconnect_1_dma_ftdi_usb3_csr_write,                                  --                                                      .write
			dma_ftdi_usb3_csr_read                                      => mm_interconnect_1_dma_ftdi_usb3_csr_read,                                   --                                                      .read
			dma_ftdi_usb3_csr_readdata                                  => mm_interconnect_1_dma_ftdi_usb3_csr_readdata,                               --                                                      .readdata
			dma_ftdi_usb3_csr_writedata                                 => mm_interconnect_1_dma_ftdi_usb3_csr_writedata,                              --                                                      .writedata
			dma_ftdi_usb3_csr_byteenable                                => mm_interconnect_1_dma_ftdi_usb3_csr_byteenable,                             --                                                      .byteenable
			dma_ftdi_usb3_descriptor_slave_write                        => mm_interconnect_1_dma_ftdi_usb3_descriptor_slave_write,                     --                        dma_ftdi_usb3_descriptor_slave.write
			dma_ftdi_usb3_descriptor_slave_writedata                    => mm_interconnect_1_dma_ftdi_usb3_descriptor_slave_writedata,                 --                                                      .writedata
			dma_ftdi_usb3_descriptor_slave_byteenable                   => mm_interconnect_1_dma_ftdi_usb3_descriptor_slave_byteenable,                --                                                      .byteenable
			dma_ftdi_usb3_descriptor_slave_waitrequest                  => mm_interconnect_1_dma_ftdi_usb3_descriptor_slave_waitrequest,               --                                                      .waitrequest
			ext_flash_uas_address                                       => mm_interconnect_1_ext_flash_uas_address,                                    --                                         ext_flash_uas.address
			ext_flash_uas_write                                         => mm_interconnect_1_ext_flash_uas_write,                                      --                                                      .write
			ext_flash_uas_read                                          => mm_interconnect_1_ext_flash_uas_read,                                       --                                                      .read
			ext_flash_uas_readdata                                      => mm_interconnect_1_ext_flash_uas_readdata,                                   --                                                      .readdata
			ext_flash_uas_writedata                                     => mm_interconnect_1_ext_flash_uas_writedata,                                  --                                                      .writedata
			ext_flash_uas_burstcount                                    => mm_interconnect_1_ext_flash_uas_burstcount,                                 --                                                      .burstcount
			ext_flash_uas_byteenable                                    => mm_interconnect_1_ext_flash_uas_byteenable,                                 --                                                      .byteenable
			ext_flash_uas_readdatavalid                                 => mm_interconnect_1_ext_flash_uas_readdatavalid,                              --                                                      .readdatavalid
			ext_flash_uas_waitrequest                                   => mm_interconnect_1_ext_flash_uas_waitrequest,                                --                                                      .waitrequest
			ext_flash_uas_lock                                          => mm_interconnect_1_ext_flash_uas_lock,                                       --                                                      .lock
			ext_flash_uas_debugaccess                                   => mm_interconnect_1_ext_flash_uas_debugaccess,                                --                                                      .debugaccess
			FTDI_USB3_0_avalon_slave_config_address                     => mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_address,                  --                       FTDI_USB3_0_avalon_slave_config.address
			FTDI_USB3_0_avalon_slave_config_write                       => mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_write,                    --                                                      .write
			FTDI_USB3_0_avalon_slave_config_read                        => mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_read,                     --                                                      .read
			FTDI_USB3_0_avalon_slave_config_readdata                    => mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_readdata,                 --                                                      .readdata
			FTDI_USB3_0_avalon_slave_config_writedata                   => mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_writedata,                --                                                      .writedata
			FTDI_USB3_0_avalon_slave_config_byteenable                  => mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_byteenable,               --                                                      .byteenable
			FTDI_USB3_0_avalon_slave_config_waitrequest                 => mm_interconnect_1_ftdi_usb3_0_avalon_slave_config_waitrequest,              --                                                      .waitrequest
			jtag_uart_0_avalon_jtag_slave_address                       => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address,                    --                         jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                         => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write,                      --                                                      .write
			jtag_uart_0_avalon_jtag_slave_read                          => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read,                       --                                                      .read
			jtag_uart_0_avalon_jtag_slave_readdata                      => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata,                   --                                                      .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                     => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata,                  --                                                      .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                   => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest,                --                                                      .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                    => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect,                 --                                                      .chipselect
			nios2_gen2_0_debug_mem_slave_address                        => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address,                     --                          nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                          => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write,                       --                                                      .write
			nios2_gen2_0_debug_mem_slave_read                           => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read,                        --                                                      .read
			nios2_gen2_0_debug_mem_slave_readdata                       => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata,                    --                                                      .readdata
			nios2_gen2_0_debug_mem_slave_writedata                      => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata,                   --                                                      .writedata
			nios2_gen2_0_debug_mem_slave_byteenable                     => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable,                  --                                                      .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                    => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest,                 --                                                      .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                    => mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess,                 --                                                      .debugaccess
			onchip_memory_s1_address                                    => mm_interconnect_1_onchip_memory_s1_address,                                 --                                      onchip_memory_s1.address
			onchip_memory_s1_write                                      => mm_interconnect_1_onchip_memory_s1_write,                                   --                                                      .write
			onchip_memory_s1_readdata                                   => mm_interconnect_1_onchip_memory_s1_readdata,                                --                                                      .readdata
			onchip_memory_s1_writedata                                  => mm_interconnect_1_onchip_memory_s1_writedata,                               --                                                      .writedata
			onchip_memory_s1_byteenable                                 => mm_interconnect_1_onchip_memory_s1_byteenable,                              --                                                      .byteenable
			onchip_memory_s1_chipselect                                 => mm_interconnect_1_onchip_memory_s1_chipselect,                              --                                                      .chipselect
			onchip_memory_s1_clken                                      => mm_interconnect_1_onchip_memory_s1_clken,                                   --                                                      .clken
			rmap_mem_nfee_comm_1_avalon_rmap_slave_0_address            => mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_address,         --              rmap_mem_nfee_comm_1_avalon_rmap_slave_0.address
			rmap_mem_nfee_comm_1_avalon_rmap_slave_0_write              => mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_write,           --                                                      .write
			rmap_mem_nfee_comm_1_avalon_rmap_slave_0_read               => mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_read,            --                                                      .read
			rmap_mem_nfee_comm_1_avalon_rmap_slave_0_readdata           => mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_readdata,        --                                                      .readdata
			rmap_mem_nfee_comm_1_avalon_rmap_slave_0_writedata          => mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_writedata,       --                                                      .writedata
			rmap_mem_nfee_comm_1_avalon_rmap_slave_0_byteenable         => mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_byteenable,      --                                                      .byteenable
			rmap_mem_nfee_comm_1_avalon_rmap_slave_0_waitrequest        => mm_interconnect_1_rmap_mem_nfee_comm_1_avalon_rmap_slave_0_waitrequest,     --                                                      .waitrequest
			rmap_mem_nfee_comm_2_avalon_rmap_slave_0_address            => mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_address,         --              rmap_mem_nfee_comm_2_avalon_rmap_slave_0.address
			rmap_mem_nfee_comm_2_avalon_rmap_slave_0_write              => mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_write,           --                                                      .write
			rmap_mem_nfee_comm_2_avalon_rmap_slave_0_read               => mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_read,            --                                                      .read
			rmap_mem_nfee_comm_2_avalon_rmap_slave_0_readdata           => mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_readdata,        --                                                      .readdata
			rmap_mem_nfee_comm_2_avalon_rmap_slave_0_writedata          => mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_writedata,       --                                                      .writedata
			rmap_mem_nfee_comm_2_avalon_rmap_slave_0_byteenable         => mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_byteenable,      --                                                      .byteenable
			rmap_mem_nfee_comm_2_avalon_rmap_slave_0_waitrequest        => mm_interconnect_1_rmap_mem_nfee_comm_2_avalon_rmap_slave_0_waitrequest,     --                                                      .waitrequest
			rmap_mem_nfee_comm_3_avalon_rmap_slave_0_address            => mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_address,         --              rmap_mem_nfee_comm_3_avalon_rmap_slave_0.address
			rmap_mem_nfee_comm_3_avalon_rmap_slave_0_write              => mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_write,           --                                                      .write
			rmap_mem_nfee_comm_3_avalon_rmap_slave_0_read               => mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_read,            --                                                      .read
			rmap_mem_nfee_comm_3_avalon_rmap_slave_0_readdata           => mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_readdata,        --                                                      .readdata
			rmap_mem_nfee_comm_3_avalon_rmap_slave_0_writedata          => mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_writedata,       --                                                      .writedata
			rmap_mem_nfee_comm_3_avalon_rmap_slave_0_byteenable         => mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_byteenable,      --                                                      .byteenable
			rmap_mem_nfee_comm_3_avalon_rmap_slave_0_waitrequest        => mm_interconnect_1_rmap_mem_nfee_comm_3_avalon_rmap_slave_0_waitrequest,     --                                                      .waitrequest
			rmap_mem_nfee_comm_4_avalon_rmap_slave_0_address            => mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_address,         --              rmap_mem_nfee_comm_4_avalon_rmap_slave_0.address
			rmap_mem_nfee_comm_4_avalon_rmap_slave_0_write              => mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_write,           --                                                      .write
			rmap_mem_nfee_comm_4_avalon_rmap_slave_0_read               => mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_read,            --                                                      .read
			rmap_mem_nfee_comm_4_avalon_rmap_slave_0_readdata           => mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_readdata,        --                                                      .readdata
			rmap_mem_nfee_comm_4_avalon_rmap_slave_0_writedata          => mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_writedata,       --                                                      .writedata
			rmap_mem_nfee_comm_4_avalon_rmap_slave_0_byteenable         => mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_byteenable,      --                                                      .byteenable
			rmap_mem_nfee_comm_4_avalon_rmap_slave_0_waitrequest        => mm_interconnect_1_rmap_mem_nfee_comm_4_avalon_rmap_slave_0_waitrequest,     --                                                      .waitrequest
			rmap_mem_nfee_comm_5_avalon_rmap_slave_0_address            => mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_address,         --              rmap_mem_nfee_comm_5_avalon_rmap_slave_0.address
			rmap_mem_nfee_comm_5_avalon_rmap_slave_0_write              => mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_write,           --                                                      .write
			rmap_mem_nfee_comm_5_avalon_rmap_slave_0_read               => mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_read,            --                                                      .read
			rmap_mem_nfee_comm_5_avalon_rmap_slave_0_readdata           => mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_readdata,        --                                                      .readdata
			rmap_mem_nfee_comm_5_avalon_rmap_slave_0_writedata          => mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_writedata,       --                                                      .writedata
			rmap_mem_nfee_comm_5_avalon_rmap_slave_0_byteenable         => mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_byteenable,      --                                                      .byteenable
			rmap_mem_nfee_comm_5_avalon_rmap_slave_0_waitrequest        => mm_interconnect_1_rmap_mem_nfee_comm_5_avalon_rmap_slave_0_waitrequest,     --                                                      .waitrequest
			rmap_mem_nfee_comm_6_avalon_rmap_slave_0_address            => mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_address,         --              rmap_mem_nfee_comm_6_avalon_rmap_slave_0.address
			rmap_mem_nfee_comm_6_avalon_rmap_slave_0_write              => mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_write,           --                                                      .write
			rmap_mem_nfee_comm_6_avalon_rmap_slave_0_read               => mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_read,            --                                                      .read
			rmap_mem_nfee_comm_6_avalon_rmap_slave_0_readdata           => mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_readdata,        --                                                      .readdata
			rmap_mem_nfee_comm_6_avalon_rmap_slave_0_writedata          => mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_writedata,       --                                                      .writedata
			rmap_mem_nfee_comm_6_avalon_rmap_slave_0_byteenable         => mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_byteenable,      --                                                      .byteenable
			rmap_mem_nfee_comm_6_avalon_rmap_slave_0_waitrequest        => mm_interconnect_1_rmap_mem_nfee_comm_6_avalon_rmap_slave_0_waitrequest,     --                                                      .waitrequest
			sysid_qsys_control_slave_address                            => mm_interconnect_1_sysid_qsys_control_slave_address,                         --                              sysid_qsys_control_slave.address
			sysid_qsys_control_slave_readdata                           => mm_interconnect_1_sysid_qsys_control_slave_readdata                         --                                                      .readdata
		);

	mm_interconnect_2 : component MebX_Qsys_Project_mm_interconnect_2
		port map (
			clk_50_clk_clk                                                         => clk50_clk,                                                                              --                                                       clk_50_clk.clk
			Altera_UP_SD_Card_Avalon_Interface_0_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                                                     -- Altera_UP_SD_Card_Avalon_Interface_0_reset_reset_bridge_in_reset.reset
			clock_bridge_afi_50_m0_reset_reset_bridge_in_reset_reset               => rst_controller_009_reset_out_reset,                                                     --               clock_bridge_afi_50_m0_reset_reset_bridge_in_reset.reset
			rs232_uart_reset_reset_bridge_in_reset_reset                           => rst_controller_013_reset_out_reset,                                                     --                           rs232_uart_reset_reset_bridge_in_reset.reset
			sync_reset_reset_bridge_in_reset_reset                                 => rst_controller_014_reset_out_reset,                                                     --                                 sync_reset_reset_bridge_in_reset.reset
			clock_bridge_afi_50_m0_address                                         => clock_bridge_afi_50_m0_address,                                                         --                                           clock_bridge_afi_50_m0.address
			clock_bridge_afi_50_m0_waitrequest                                     => clock_bridge_afi_50_m0_waitrequest,                                                     --                                                                 .waitrequest
			clock_bridge_afi_50_m0_burstcount                                      => clock_bridge_afi_50_m0_burstcount,                                                      --                                                                 .burstcount
			clock_bridge_afi_50_m0_byteenable                                      => clock_bridge_afi_50_m0_byteenable,                                                      --                                                                 .byteenable
			clock_bridge_afi_50_m0_read                                            => clock_bridge_afi_50_m0_read,                                                            --                                                                 .read
			clock_bridge_afi_50_m0_readdata                                        => clock_bridge_afi_50_m0_readdata,                                                        --                                                                 .readdata
			clock_bridge_afi_50_m0_readdatavalid                                   => clock_bridge_afi_50_m0_readdatavalid,                                                   --                                                                 .readdatavalid
			clock_bridge_afi_50_m0_write                                           => clock_bridge_afi_50_m0_write,                                                           --                                                                 .write
			clock_bridge_afi_50_m0_writedata                                       => clock_bridge_afi_50_m0_writedata,                                                       --                                                                 .writedata
			clock_bridge_afi_50_m0_debugaccess                                     => clock_bridge_afi_50_m0_debugaccess,                                                     --                                                                 .debugaccess
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_address       => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_address,     --         Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave.address
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_write         => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_write,       --                                                                 .write
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_read          => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_read,        --                                                                 .read
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_readdata      => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_readdata,    --                                                                 .readdata
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_writedata     => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_writedata,   --                                                                 .writedata
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_byteenable    => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_byteenable,  --                                                                 .byteenable
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_waitrequest   => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_waitrequest, --                                                                 .waitrequest
			Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_chipselect    => mm_interconnect_2_altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_chipselect,  --                                                                 .chipselect
			csense_adc_fo_s1_address                                               => mm_interconnect_2_csense_adc_fo_s1_address,                                             --                                                 csense_adc_fo_s1.address
			csense_adc_fo_s1_write                                                 => mm_interconnect_2_csense_adc_fo_s1_write,                                               --                                                                 .write
			csense_adc_fo_s1_readdata                                              => mm_interconnect_2_csense_adc_fo_s1_readdata,                                            --                                                                 .readdata
			csense_adc_fo_s1_writedata                                             => mm_interconnect_2_csense_adc_fo_s1_writedata,                                           --                                                                 .writedata
			csense_adc_fo_s1_chipselect                                            => mm_interconnect_2_csense_adc_fo_s1_chipselect,                                          --                                                                 .chipselect
			csense_cs_n_s1_address                                                 => mm_interconnect_2_csense_cs_n_s1_address,                                               --                                                   csense_cs_n_s1.address
			csense_cs_n_s1_write                                                   => mm_interconnect_2_csense_cs_n_s1_write,                                                 --                                                                 .write
			csense_cs_n_s1_readdata                                                => mm_interconnect_2_csense_cs_n_s1_readdata,                                              --                                                                 .readdata
			csense_cs_n_s1_writedata                                               => mm_interconnect_2_csense_cs_n_s1_writedata,                                             --                                                                 .writedata
			csense_cs_n_s1_chipselect                                              => mm_interconnect_2_csense_cs_n_s1_chipselect,                                            --                                                                 .chipselect
			csense_sck_s1_address                                                  => mm_interconnect_2_csense_sck_s1_address,                                                --                                                    csense_sck_s1.address
			csense_sck_s1_write                                                    => mm_interconnect_2_csense_sck_s1_write,                                                  --                                                                 .write
			csense_sck_s1_readdata                                                 => mm_interconnect_2_csense_sck_s1_readdata,                                               --                                                                 .readdata
			csense_sck_s1_writedata                                                => mm_interconnect_2_csense_sck_s1_writedata,                                              --                                                                 .writedata
			csense_sck_s1_chipselect                                               => mm_interconnect_2_csense_sck_s1_chipselect,                                             --                                                                 .chipselect
			csense_sdi_s1_address                                                  => mm_interconnect_2_csense_sdi_s1_address,                                                --                                                    csense_sdi_s1.address
			csense_sdi_s1_write                                                    => mm_interconnect_2_csense_sdi_s1_write,                                                  --                                                                 .write
			csense_sdi_s1_readdata                                                 => mm_interconnect_2_csense_sdi_s1_readdata,                                               --                                                                 .readdata
			csense_sdi_s1_writedata                                                => mm_interconnect_2_csense_sdi_s1_writedata,                                              --                                                                 .writedata
			csense_sdi_s1_chipselect                                               => mm_interconnect_2_csense_sdi_s1_chipselect,                                             --                                                                 .chipselect
			csense_sdo_s1_address                                                  => mm_interconnect_2_csense_sdo_s1_address,                                                --                                                    csense_sdo_s1.address
			csense_sdo_s1_readdata                                                 => mm_interconnect_2_csense_sdo_s1_readdata,                                               --                                                                 .readdata
			m1_ddr2_i2c_scl_s1_address                                             => mm_interconnect_2_m1_ddr2_i2c_scl_s1_address,                                           --                                               m1_ddr2_i2c_scl_s1.address
			m1_ddr2_i2c_scl_s1_write                                               => mm_interconnect_2_m1_ddr2_i2c_scl_s1_write,                                             --                                                                 .write
			m1_ddr2_i2c_scl_s1_readdata                                            => mm_interconnect_2_m1_ddr2_i2c_scl_s1_readdata,                                          --                                                                 .readdata
			m1_ddr2_i2c_scl_s1_writedata                                           => mm_interconnect_2_m1_ddr2_i2c_scl_s1_writedata,                                         --                                                                 .writedata
			m1_ddr2_i2c_scl_s1_chipselect                                          => mm_interconnect_2_m1_ddr2_i2c_scl_s1_chipselect,                                        --                                                                 .chipselect
			m1_ddr2_i2c_sda_s1_address                                             => mm_interconnect_2_m1_ddr2_i2c_sda_s1_address,                                           --                                               m1_ddr2_i2c_sda_s1.address
			m1_ddr2_i2c_sda_s1_write                                               => mm_interconnect_2_m1_ddr2_i2c_sda_s1_write,                                             --                                                                 .write
			m1_ddr2_i2c_sda_s1_readdata                                            => mm_interconnect_2_m1_ddr2_i2c_sda_s1_readdata,                                          --                                                                 .readdata
			m1_ddr2_i2c_sda_s1_writedata                                           => mm_interconnect_2_m1_ddr2_i2c_sda_s1_writedata,                                         --                                                                 .writedata
			m1_ddr2_i2c_sda_s1_chipselect                                          => mm_interconnect_2_m1_ddr2_i2c_sda_s1_chipselect,                                        --                                                                 .chipselect
			m2_ddr2_i2c_scl_s1_address                                             => mm_interconnect_2_m2_ddr2_i2c_scl_s1_address,                                           --                                               m2_ddr2_i2c_scl_s1.address
			m2_ddr2_i2c_scl_s1_write                                               => mm_interconnect_2_m2_ddr2_i2c_scl_s1_write,                                             --                                                                 .write
			m2_ddr2_i2c_scl_s1_readdata                                            => mm_interconnect_2_m2_ddr2_i2c_scl_s1_readdata,                                          --                                                                 .readdata
			m2_ddr2_i2c_scl_s1_writedata                                           => mm_interconnect_2_m2_ddr2_i2c_scl_s1_writedata,                                         --                                                                 .writedata
			m2_ddr2_i2c_scl_s1_chipselect                                          => mm_interconnect_2_m2_ddr2_i2c_scl_s1_chipselect,                                        --                                                                 .chipselect
			m2_ddr2_i2c_sda_s1_address                                             => mm_interconnect_2_m2_ddr2_i2c_sda_s1_address,                                           --                                               m2_ddr2_i2c_sda_s1.address
			m2_ddr2_i2c_sda_s1_write                                               => mm_interconnect_2_m2_ddr2_i2c_sda_s1_write,                                             --                                                                 .write
			m2_ddr2_i2c_sda_s1_readdata                                            => mm_interconnect_2_m2_ddr2_i2c_sda_s1_readdata,                                          --                                                                 .readdata
			m2_ddr2_i2c_sda_s1_writedata                                           => mm_interconnect_2_m2_ddr2_i2c_sda_s1_writedata,                                         --                                                                 .writedata
			m2_ddr2_i2c_sda_s1_chipselect                                          => mm_interconnect_2_m2_ddr2_i2c_sda_s1_chipselect,                                        --                                                                 .chipselect
			pio_BUTTON_s1_address                                                  => mm_interconnect_2_pio_button_s1_address,                                                --                                                    pio_BUTTON_s1.address
			pio_BUTTON_s1_readdata                                                 => mm_interconnect_2_pio_button_s1_readdata,                                               --                                                                 .readdata
			pio_ctrl_io_lvds_s1_address                                            => mm_interconnect_2_pio_ctrl_io_lvds_s1_address,                                          --                                              pio_ctrl_io_lvds_s1.address
			pio_ctrl_io_lvds_s1_write                                              => mm_interconnect_2_pio_ctrl_io_lvds_s1_write,                                            --                                                                 .write
			pio_ctrl_io_lvds_s1_readdata                                           => mm_interconnect_2_pio_ctrl_io_lvds_s1_readdata,                                         --                                                                 .readdata
			pio_ctrl_io_lvds_s1_writedata                                          => mm_interconnect_2_pio_ctrl_io_lvds_s1_writedata,                                        --                                                                 .writedata
			pio_ctrl_io_lvds_s1_chipselect                                         => mm_interconnect_2_pio_ctrl_io_lvds_s1_chipselect,                                       --                                                                 .chipselect
			pio_DIP_s1_address                                                     => mm_interconnect_2_pio_dip_s1_address,                                                   --                                                       pio_DIP_s1.address
			pio_DIP_s1_readdata                                                    => mm_interconnect_2_pio_dip_s1_readdata,                                                  --                                                                 .readdata
			pio_EXT_s1_address                                                     => mm_interconnect_2_pio_ext_s1_address,                                                   --                                                       pio_EXT_s1.address
			pio_EXT_s1_readdata                                                    => mm_interconnect_2_pio_ext_s1_readdata,                                                  --                                                                 .readdata
			pio_LED_s1_address                                                     => mm_interconnect_2_pio_led_s1_address,                                                   --                                                       pio_LED_s1.address
			pio_LED_s1_write                                                       => mm_interconnect_2_pio_led_s1_write,                                                     --                                                                 .write
			pio_LED_s1_readdata                                                    => mm_interconnect_2_pio_led_s1_readdata,                                                  --                                                                 .readdata
			pio_LED_s1_writedata                                                   => mm_interconnect_2_pio_led_s1_writedata,                                                 --                                                                 .writedata
			pio_LED_s1_chipselect                                                  => mm_interconnect_2_pio_led_s1_chipselect,                                                --                                                                 .chipselect
			pio_LED_painel_s1_address                                              => mm_interconnect_2_pio_led_painel_s1_address,                                            --                                                pio_LED_painel_s1.address
			pio_LED_painel_s1_write                                                => mm_interconnect_2_pio_led_painel_s1_write,                                              --                                                                 .write
			pio_LED_painel_s1_readdata                                             => mm_interconnect_2_pio_led_painel_s1_readdata,                                           --                                                                 .readdata
			pio_LED_painel_s1_writedata                                            => mm_interconnect_2_pio_led_painel_s1_writedata,                                          --                                                                 .writedata
			pio_LED_painel_s1_chipselect                                           => mm_interconnect_2_pio_led_painel_s1_chipselect,                                         --                                                                 .chipselect
			rs232_uart_s1_address                                                  => mm_interconnect_2_rs232_uart_s1_address,                                                --                                                    rs232_uart_s1.address
			rs232_uart_s1_write                                                    => mm_interconnect_2_rs232_uart_s1_write,                                                  --                                                                 .write
			rs232_uart_s1_read                                                     => mm_interconnect_2_rs232_uart_s1_read,                                                   --                                                                 .read
			rs232_uart_s1_readdata                                                 => mm_interconnect_2_rs232_uart_s1_readdata,                                               --                                                                 .readdata
			rs232_uart_s1_writedata                                                => mm_interconnect_2_rs232_uart_s1_writedata,                                              --                                                                 .writedata
			rs232_uart_s1_begintransfer                                            => mm_interconnect_2_rs232_uart_s1_begintransfer,                                          --                                                                 .begintransfer
			rs232_uart_s1_chipselect                                               => mm_interconnect_2_rs232_uart_s1_chipselect,                                             --                                                                 .chipselect
			rst_controller_avalon_rst_controller_slave_address                     => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_address,                   --                       rst_controller_avalon_rst_controller_slave.address
			rst_controller_avalon_rst_controller_slave_write                       => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_write,                     --                                                                 .write
			rst_controller_avalon_rst_controller_slave_read                        => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_read,                      --                                                                 .read
			rst_controller_avalon_rst_controller_slave_readdata                    => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_readdata,                  --                                                                 .readdata
			rst_controller_avalon_rst_controller_slave_writedata                   => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_writedata,                 --                                                                 .writedata
			rst_controller_avalon_rst_controller_slave_waitrequest                 => mm_interconnect_2_rst_controller_avalon_rst_controller_slave_waitrequest,               --                                                                 .waitrequest
			rtcc_alarm_s1_address                                                  => mm_interconnect_2_rtcc_alarm_s1_address,                                                --                                                    rtcc_alarm_s1.address
			rtcc_alarm_s1_readdata                                                 => mm_interconnect_2_rtcc_alarm_s1_readdata,                                               --                                                                 .readdata
			rtcc_cs_n_s1_address                                                   => mm_interconnect_2_rtcc_cs_n_s1_address,                                                 --                                                     rtcc_cs_n_s1.address
			rtcc_cs_n_s1_write                                                     => mm_interconnect_2_rtcc_cs_n_s1_write,                                                   --                                                                 .write
			rtcc_cs_n_s1_readdata                                                  => mm_interconnect_2_rtcc_cs_n_s1_readdata,                                                --                                                                 .readdata
			rtcc_cs_n_s1_writedata                                                 => mm_interconnect_2_rtcc_cs_n_s1_writedata,                                               --                                                                 .writedata
			rtcc_cs_n_s1_chipselect                                                => mm_interconnect_2_rtcc_cs_n_s1_chipselect,                                              --                                                                 .chipselect
			rtcc_sck_s1_address                                                    => mm_interconnect_2_rtcc_sck_s1_address,                                                  --                                                      rtcc_sck_s1.address
			rtcc_sck_s1_write                                                      => mm_interconnect_2_rtcc_sck_s1_write,                                                    --                                                                 .write
			rtcc_sck_s1_readdata                                                   => mm_interconnect_2_rtcc_sck_s1_readdata,                                                 --                                                                 .readdata
			rtcc_sck_s1_writedata                                                  => mm_interconnect_2_rtcc_sck_s1_writedata,                                                --                                                                 .writedata
			rtcc_sck_s1_chipselect                                                 => mm_interconnect_2_rtcc_sck_s1_chipselect,                                               --                                                                 .chipselect
			rtcc_sdi_s1_address                                                    => mm_interconnect_2_rtcc_sdi_s1_address,                                                  --                                                      rtcc_sdi_s1.address
			rtcc_sdi_s1_write                                                      => mm_interconnect_2_rtcc_sdi_s1_write,                                                    --                                                                 .write
			rtcc_sdi_s1_readdata                                                   => mm_interconnect_2_rtcc_sdi_s1_readdata,                                                 --                                                                 .readdata
			rtcc_sdi_s1_writedata                                                  => mm_interconnect_2_rtcc_sdi_s1_writedata,                                                --                                                                 .writedata
			rtcc_sdi_s1_chipselect                                                 => mm_interconnect_2_rtcc_sdi_s1_chipselect,                                               --                                                                 .chipselect
			rtcc_sdo_s1_address                                                    => mm_interconnect_2_rtcc_sdo_s1_address,                                                  --                                                      rtcc_sdo_s1.address
			rtcc_sdo_s1_readdata                                                   => mm_interconnect_2_rtcc_sdo_s1_readdata,                                                 --                                                                 .readdata
			sd_card_wp_n_s1_address                                                => mm_interconnect_2_sd_card_wp_n_s1_address,                                              --                                                  sd_card_wp_n_s1.address
			sd_card_wp_n_s1_readdata                                               => mm_interconnect_2_sd_card_wp_n_s1_readdata,                                             --                                                                 .readdata
			SEVEN_SEGMENT_CONTROLLER_0_SSDP_avalon_slave_address                   => mm_interconnect_2_seven_segment_controller_0_ssdp_avalon_slave_address,                 --                     SEVEN_SEGMENT_CONTROLLER_0_SSDP_avalon_slave.address
			SEVEN_SEGMENT_CONTROLLER_0_SSDP_avalon_slave_write                     => mm_interconnect_2_seven_segment_controller_0_ssdp_avalon_slave_write,                   --                                                                 .write
			SEVEN_SEGMENT_CONTROLLER_0_SSDP_avalon_slave_writedata                 => mm_interconnect_2_seven_segment_controller_0_ssdp_avalon_slave_writedata,               --                                                                 .writedata
			sync_avalon_mm_slave_address                                           => mm_interconnect_2_sync_avalon_mm_slave_address,                                         --                                             sync_avalon_mm_slave.address
			sync_avalon_mm_slave_write                                             => mm_interconnect_2_sync_avalon_mm_slave_write,                                           --                                                                 .write
			sync_avalon_mm_slave_read                                              => mm_interconnect_2_sync_avalon_mm_slave_read,                                            --                                                                 .read
			sync_avalon_mm_slave_readdata                                          => mm_interconnect_2_sync_avalon_mm_slave_readdata,                                        --                                                                 .readdata
			sync_avalon_mm_slave_writedata                                         => mm_interconnect_2_sync_avalon_mm_slave_writedata,                                       --                                                                 .writedata
			sync_avalon_mm_slave_byteenable                                        => mm_interconnect_2_sync_avalon_mm_slave_byteenable,                                      --                                                                 .byteenable
			sync_avalon_mm_slave_waitrequest                                       => mm_interconnect_2_sync_avalon_mm_slave_waitrequest,                                     --                                                                 .waitrequest
			temp_scl_s1_address                                                    => mm_interconnect_2_temp_scl_s1_address,                                                  --                                                      temp_scl_s1.address
			temp_scl_s1_write                                                      => mm_interconnect_2_temp_scl_s1_write,                                                    --                                                                 .write
			temp_scl_s1_readdata                                                   => mm_interconnect_2_temp_scl_s1_readdata,                                                 --                                                                 .readdata
			temp_scl_s1_writedata                                                  => mm_interconnect_2_temp_scl_s1_writedata,                                                --                                                                 .writedata
			temp_scl_s1_chipselect                                                 => mm_interconnect_2_temp_scl_s1_chipselect,                                               --                                                                 .chipselect
			temp_sda_s1_address                                                    => mm_interconnect_2_temp_sda_s1_address,                                                  --                                                      temp_sda_s1.address
			temp_sda_s1_write                                                      => mm_interconnect_2_temp_sda_s1_write,                                                    --                                                                 .write
			temp_sda_s1_readdata                                                   => mm_interconnect_2_temp_sda_s1_readdata,                                                 --                                                                 .readdata
			temp_sda_s1_writedata                                                  => mm_interconnect_2_temp_sda_s1_writedata,                                                --                                                                 .writedata
			temp_sda_s1_chipselect                                                 => mm_interconnect_2_temp_sda_s1_chipselect,                                               --                                                                 .chipselect
			timer_1ms_s1_address                                                   => mm_interconnect_2_timer_1ms_s1_address,                                                 --                                                     timer_1ms_s1.address
			timer_1ms_s1_write                                                     => mm_interconnect_2_timer_1ms_s1_write,                                                   --                                                                 .write
			timer_1ms_s1_readdata                                                  => mm_interconnect_2_timer_1ms_s1_readdata,                                                --                                                                 .readdata
			timer_1ms_s1_writedata                                                 => mm_interconnect_2_timer_1ms_s1_writedata,                                               --                                                                 .writedata
			timer_1ms_s1_chipselect                                                => mm_interconnect_2_timer_1ms_s1_chipselect,                                              --                                                                 .chipselect
			timer_1us_s1_address                                                   => mm_interconnect_2_timer_1us_s1_address,                                                 --                                                     timer_1us_s1.address
			timer_1us_s1_write                                                     => mm_interconnect_2_timer_1us_s1_write,                                                   --                                                                 .write
			timer_1us_s1_readdata                                                  => mm_interconnect_2_timer_1us_s1_readdata,                                                --                                                                 .readdata
			timer_1us_s1_writedata                                                 => mm_interconnect_2_timer_1us_s1_writedata,                                               --                                                                 .writedata
			timer_1us_s1_chipselect                                                => mm_interconnect_2_timer_1us_s1_chipselect                                               --                                                                 .chipselect
		);

	mm_interconnect_3 : component MebX_Qsys_Project_mm_interconnect_3
		port map (
			m1_ddr2_memory_afi_clk_clk                                      => m1_ddr2_memory_afi_clk_clk,                              --                                    m1_ddr2_memory_afi_clk.clk
			m1_ddr2_memory_afi_half_clk_clk                                 => m1_ddr2_memory_afi_half_clk_clk,                         --                               m1_ddr2_memory_afi_half_clk.clk
			m1_clock_bridge_m0_reset_reset_bridge_in_reset_reset            => rst_controller_011_reset_out_reset,                      --            m1_clock_bridge_m0_reset_reset_bridge_in_reset.reset
			m1_ddr2_memory_avl_translator_reset_reset_bridge_in_reset_reset => rst_controller_016_reset_out_reset,                      -- m1_ddr2_memory_avl_translator_reset_reset_bridge_in_reset.reset
			m1_ddr2_memory_soft_reset_reset_bridge_in_reset_reset           => rst_controller_016_reset_out_reset,                      --           m1_ddr2_memory_soft_reset_reset_bridge_in_reset.reset
			m1_clock_bridge_m0_address                                      => m1_clock_bridge_m0_address,                              --                                        m1_clock_bridge_m0.address
			m1_clock_bridge_m0_waitrequest                                  => m1_clock_bridge_m0_waitrequest,                          --                                                          .waitrequest
			m1_clock_bridge_m0_burstcount                                   => m1_clock_bridge_m0_burstcount,                           --                                                          .burstcount
			m1_clock_bridge_m0_byteenable                                   => m1_clock_bridge_m0_byteenable,                           --                                                          .byteenable
			m1_clock_bridge_m0_read                                         => m1_clock_bridge_m0_read,                                 --                                                          .read
			m1_clock_bridge_m0_readdata                                     => m1_clock_bridge_m0_readdata,                             --                                                          .readdata
			m1_clock_bridge_m0_readdatavalid                                => m1_clock_bridge_m0_readdatavalid,                        --                                                          .readdatavalid
			m1_clock_bridge_m0_write                                        => m1_clock_bridge_m0_write,                                --                                                          .write
			m1_clock_bridge_m0_writedata                                    => m1_clock_bridge_m0_writedata,                            --                                                          .writedata
			m1_clock_bridge_m0_debugaccess                                  => m1_clock_bridge_m0_debugaccess,                          --                                                          .debugaccess
			m1_ddr2_memory_avl_address                                      => mm_interconnect_3_m1_ddr2_memory_avl_address,            --                                        m1_ddr2_memory_avl.address
			m1_ddr2_memory_avl_write                                        => mm_interconnect_3_m1_ddr2_memory_avl_write,              --                                                          .write
			m1_ddr2_memory_avl_read                                         => mm_interconnect_3_m1_ddr2_memory_avl_read,               --                                                          .read
			m1_ddr2_memory_avl_readdata                                     => mm_interconnect_3_m1_ddr2_memory_avl_readdata,           --                                                          .readdata
			m1_ddr2_memory_avl_writedata                                    => mm_interconnect_3_m1_ddr2_memory_avl_writedata,          --                                                          .writedata
			m1_ddr2_memory_avl_beginbursttransfer                           => mm_interconnect_3_m1_ddr2_memory_avl_beginbursttransfer, --                                                          .beginbursttransfer
			m1_ddr2_memory_avl_burstcount                                   => mm_interconnect_3_m1_ddr2_memory_avl_burstcount,         --                                                          .burstcount
			m1_ddr2_memory_avl_byteenable                                   => mm_interconnect_3_m1_ddr2_memory_avl_byteenable,         --                                                          .byteenable
			m1_ddr2_memory_avl_readdatavalid                                => mm_interconnect_3_m1_ddr2_memory_avl_readdatavalid,      --                                                          .readdatavalid
			m1_ddr2_memory_avl_waitrequest                                  => mm_interconnect_3_m1_ddr2_memory_avl_inv                 --                                                          .waitrequest
		);

	mm_interconnect_4 : component MebX_Qsys_Project_mm_interconnect_4
		port map (
			clk_100_clk_clk                                   => m2_ddr2_memory_afi_half_clk_clk,                             --                                 clk_100_clk.clk
			dma_ftdi_usb3_reset_n_reset_bridge_in_reset_reset => rst_controller_008_reset_out_reset,                          -- dma_ftdi_usb3_reset_n_reset_bridge_in_reset.reset
			dma_ftdi_usb3_mm_read_address                     => dma_ftdi_usb3_mm_read_address,                               --                       dma_ftdi_usb3_mm_read.address
			dma_ftdi_usb3_mm_read_waitrequest                 => dma_ftdi_usb3_mm_read_waitrequest,                           --                                            .waitrequest
			dma_ftdi_usb3_mm_read_byteenable                  => dma_ftdi_usb3_mm_read_byteenable,                            --                                            .byteenable
			dma_ftdi_usb3_mm_read_read                        => dma_ftdi_usb3_mm_read_read,                                  --                                            .read
			dma_ftdi_usb3_mm_read_readdata                    => dma_ftdi_usb3_mm_read_readdata,                              --                                            .readdata
			dma_ftdi_usb3_mm_read_readdatavalid               => dma_ftdi_usb3_mm_read_readdatavalid,                         --                                            .readdatavalid
			FTDI_USB3_0_avalon_slave_data_address             => mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_address,     --               FTDI_USB3_0_avalon_slave_data.address
			FTDI_USB3_0_avalon_slave_data_write               => mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_write,       --                                            .write
			FTDI_USB3_0_avalon_slave_data_read                => mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_read,        --                                            .read
			FTDI_USB3_0_avalon_slave_data_readdata            => mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_readdata,    --                                            .readdata
			FTDI_USB3_0_avalon_slave_data_writedata           => mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_writedata,   --                                            .writedata
			FTDI_USB3_0_avalon_slave_data_waitrequest         => mm_interconnect_4_ftdi_usb3_0_avalon_slave_data_waitrequest  --                                            .waitrequest
		);

	mm_interconnect_5 : component MebX_Qsys_Project_mm_interconnect_5
		port map (
			clk_100_clk_clk                                              => m2_ddr2_memory_afi_half_clk_clk,                                           --                                            clk_100_clk.clk
			COMM_Pedreiro_v1_01_A_reset_sink_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                                        -- COMM_Pedreiro_v1_01_A_reset_sink_reset_bridge_in_reset.reset
			dma_comm_1_left_reset_n_reset_bridge_in_reset_reset          => rst_controller_008_reset_out_reset,                                        --          dma_comm_1_left_reset_n_reset_bridge_in_reset.reset
			dma_comm_1_left_mm_write_address                             => dma_comm_1_left_mm_write_address,                                          --                               dma_comm_1_left_mm_write.address
			dma_comm_1_left_mm_write_waitrequest                         => dma_comm_1_left_mm_write_waitrequest,                                      --                                                       .waitrequest
			dma_comm_1_left_mm_write_byteenable                          => dma_comm_1_left_mm_write_byteenable,                                       --                                                       .byteenable
			dma_comm_1_left_mm_write_write                               => dma_comm_1_left_mm_write_write,                                            --                                                       .write
			dma_comm_1_left_mm_write_writedata                           => dma_comm_1_left_mm_write_writedata,                                        --                                                       .writedata
			COMM_Pedreiro_v1_01_A_avalon_slave_L_buffer_address          => mm_interconnect_5_comm_pedreiro_v1_01_a_avalon_slave_l_buffer_address,     --            COMM_Pedreiro_v1_01_A_avalon_slave_L_buffer.address
			COMM_Pedreiro_v1_01_A_avalon_slave_L_buffer_write            => mm_interconnect_5_comm_pedreiro_v1_01_a_avalon_slave_l_buffer_write,       --                                                       .write
			COMM_Pedreiro_v1_01_A_avalon_slave_L_buffer_writedata        => mm_interconnect_5_comm_pedreiro_v1_01_a_avalon_slave_l_buffer_writedata,   --                                                       .writedata
			COMM_Pedreiro_v1_01_A_avalon_slave_L_buffer_waitrequest      => mm_interconnect_5_comm_pedreiro_v1_01_a_avalon_slave_l_buffer_waitrequest  --                                                       .waitrequest
		);

	mm_interconnect_6 : component MebX_Qsys_Project_mm_interconnect_6
		port map (
			clk_100_clk_clk                                              => m2_ddr2_memory_afi_half_clk_clk,                                           --                                            clk_100_clk.clk
			COMM_Pedreiro_v1_01_B_reset_sink_reset_bridge_in_reset_reset => rst_controller_003_reset_out_reset,                                        -- COMM_Pedreiro_v1_01_B_reset_sink_reset_bridge_in_reset.reset
			dma_comm_2_left_reset_n_reset_bridge_in_reset_reset          => rst_controller_008_reset_out_reset,                                        --          dma_comm_2_left_reset_n_reset_bridge_in_reset.reset
			dma_comm_2_left_mm_write_address                             => dma_comm_2_left_mm_write_address,                                          --                               dma_comm_2_left_mm_write.address
			dma_comm_2_left_mm_write_waitrequest                         => dma_comm_2_left_mm_write_waitrequest,                                      --                                                       .waitrequest
			dma_comm_2_left_mm_write_byteenable                          => dma_comm_2_left_mm_write_byteenable,                                       --                                                       .byteenable
			dma_comm_2_left_mm_write_write                               => dma_comm_2_left_mm_write_write,                                            --                                                       .write
			dma_comm_2_left_mm_write_writedata                           => dma_comm_2_left_mm_write_writedata,                                        --                                                       .writedata
			COMM_Pedreiro_v1_01_B_avalon_slave_L_buffer_address          => mm_interconnect_6_comm_pedreiro_v1_01_b_avalon_slave_l_buffer_address,     --            COMM_Pedreiro_v1_01_B_avalon_slave_L_buffer.address
			COMM_Pedreiro_v1_01_B_avalon_slave_L_buffer_write            => mm_interconnect_6_comm_pedreiro_v1_01_b_avalon_slave_l_buffer_write,       --                                                       .write
			COMM_Pedreiro_v1_01_B_avalon_slave_L_buffer_writedata        => mm_interconnect_6_comm_pedreiro_v1_01_b_avalon_slave_l_buffer_writedata,   --                                                       .writedata
			COMM_Pedreiro_v1_01_B_avalon_slave_L_buffer_waitrequest      => mm_interconnect_6_comm_pedreiro_v1_01_b_avalon_slave_l_buffer_waitrequest  --                                                       .waitrequest
		);

	mm_interconnect_7 : component MebX_Qsys_Project_mm_interconnect_7
		port map (
			clk_100_clk_clk                                              => m2_ddr2_memory_afi_half_clk_clk,                                           --                                            clk_100_clk.clk
			COMM_Pedreiro_v1_01_C_reset_sink_reset_bridge_in_reset_reset => rst_controller_004_reset_out_reset,                                        -- COMM_Pedreiro_v1_01_C_reset_sink_reset_bridge_in_reset.reset
			dma_comm_3_left_reset_n_reset_bridge_in_reset_reset          => rst_controller_008_reset_out_reset,                                        --          dma_comm_3_left_reset_n_reset_bridge_in_reset.reset
			dma_comm_3_left_mm_write_address                             => dma_comm_3_left_mm_write_address,                                          --                               dma_comm_3_left_mm_write.address
			dma_comm_3_left_mm_write_waitrequest                         => dma_comm_3_left_mm_write_waitrequest,                                      --                                                       .waitrequest
			dma_comm_3_left_mm_write_byteenable                          => dma_comm_3_left_mm_write_byteenable,                                       --                                                       .byteenable
			dma_comm_3_left_mm_write_write                               => dma_comm_3_left_mm_write_write,                                            --                                                       .write
			dma_comm_3_left_mm_write_writedata                           => dma_comm_3_left_mm_write_writedata,                                        --                                                       .writedata
			COMM_Pedreiro_v1_01_C_avalon_slave_L_buffer_address          => mm_interconnect_7_comm_pedreiro_v1_01_c_avalon_slave_l_buffer_address,     --            COMM_Pedreiro_v1_01_C_avalon_slave_L_buffer.address
			COMM_Pedreiro_v1_01_C_avalon_slave_L_buffer_write            => mm_interconnect_7_comm_pedreiro_v1_01_c_avalon_slave_l_buffer_write,       --                                                       .write
			COMM_Pedreiro_v1_01_C_avalon_slave_L_buffer_writedata        => mm_interconnect_7_comm_pedreiro_v1_01_c_avalon_slave_l_buffer_writedata,   --                                                       .writedata
			COMM_Pedreiro_v1_01_C_avalon_slave_L_buffer_waitrequest      => mm_interconnect_7_comm_pedreiro_v1_01_c_avalon_slave_l_buffer_waitrequest  --                                                       .waitrequest
		);

	mm_interconnect_8 : component MebX_Qsys_Project_mm_interconnect_8
		port map (
			clk_100_clk_clk                                              => m2_ddr2_memory_afi_half_clk_clk,                                           --                                            clk_100_clk.clk
			COMM_Pedreiro_v1_01_D_reset_sink_reset_bridge_in_reset_reset => rst_controller_005_reset_out_reset,                                        -- COMM_Pedreiro_v1_01_D_reset_sink_reset_bridge_in_reset.reset
			dma_comm_4_left_reset_n_reset_bridge_in_reset_reset          => rst_controller_008_reset_out_reset,                                        --          dma_comm_4_left_reset_n_reset_bridge_in_reset.reset
			dma_comm_4_left_mm_write_address                             => dma_comm_4_left_mm_write_address,                                          --                               dma_comm_4_left_mm_write.address
			dma_comm_4_left_mm_write_waitrequest                         => dma_comm_4_left_mm_write_waitrequest,                                      --                                                       .waitrequest
			dma_comm_4_left_mm_write_byteenable                          => dma_comm_4_left_mm_write_byteenable,                                       --                                                       .byteenable
			dma_comm_4_left_mm_write_write                               => dma_comm_4_left_mm_write_write,                                            --                                                       .write
			dma_comm_4_left_mm_write_writedata                           => dma_comm_4_left_mm_write_writedata,                                        --                                                       .writedata
			COMM_Pedreiro_v1_01_D_avalon_slave_L_buffer_address          => mm_interconnect_8_comm_pedreiro_v1_01_d_avalon_slave_l_buffer_address,     --            COMM_Pedreiro_v1_01_D_avalon_slave_L_buffer.address
			COMM_Pedreiro_v1_01_D_avalon_slave_L_buffer_write            => mm_interconnect_8_comm_pedreiro_v1_01_d_avalon_slave_l_buffer_write,       --                                                       .write
			COMM_Pedreiro_v1_01_D_avalon_slave_L_buffer_writedata        => mm_interconnect_8_comm_pedreiro_v1_01_d_avalon_slave_l_buffer_writedata,   --                                                       .writedata
			COMM_Pedreiro_v1_01_D_avalon_slave_L_buffer_waitrequest      => mm_interconnect_8_comm_pedreiro_v1_01_d_avalon_slave_l_buffer_waitrequest  --                                                       .waitrequest
		);

	mm_interconnect_9 : component MebX_Qsys_Project_mm_interconnect_9
		port map (
			clk_100_clk_clk                                              => m2_ddr2_memory_afi_half_clk_clk,                                           --                                            clk_100_clk.clk
			COMM_Pedreiro_v1_01_E_reset_sink_reset_bridge_in_reset_reset => rst_controller_006_reset_out_reset,                                        -- COMM_Pedreiro_v1_01_E_reset_sink_reset_bridge_in_reset.reset
			dma_comm_5_left_reset_n_reset_bridge_in_reset_reset          => rst_controller_008_reset_out_reset,                                        --          dma_comm_5_left_reset_n_reset_bridge_in_reset.reset
			dma_comm_5_left_mm_write_address                             => dma_comm_5_left_mm_write_address,                                          --                               dma_comm_5_left_mm_write.address
			dma_comm_5_left_mm_write_waitrequest                         => dma_comm_5_left_mm_write_waitrequest,                                      --                                                       .waitrequest
			dma_comm_5_left_mm_write_byteenable                          => dma_comm_5_left_mm_write_byteenable,                                       --                                                       .byteenable
			dma_comm_5_left_mm_write_write                               => dma_comm_5_left_mm_write_write,                                            --                                                       .write
			dma_comm_5_left_mm_write_writedata                           => dma_comm_5_left_mm_write_writedata,                                        --                                                       .writedata
			COMM_Pedreiro_v1_01_E_avalon_slave_L_buffer_address          => mm_interconnect_9_comm_pedreiro_v1_01_e_avalon_slave_l_buffer_address,     --            COMM_Pedreiro_v1_01_E_avalon_slave_L_buffer.address
			COMM_Pedreiro_v1_01_E_avalon_slave_L_buffer_write            => mm_interconnect_9_comm_pedreiro_v1_01_e_avalon_slave_l_buffer_write,       --                                                       .write
			COMM_Pedreiro_v1_01_E_avalon_slave_L_buffer_writedata        => mm_interconnect_9_comm_pedreiro_v1_01_e_avalon_slave_l_buffer_writedata,   --                                                       .writedata
			COMM_Pedreiro_v1_01_E_avalon_slave_L_buffer_waitrequest      => mm_interconnect_9_comm_pedreiro_v1_01_e_avalon_slave_l_buffer_waitrequest  --                                                       .waitrequest
		);

	mm_interconnect_10 : component MebX_Qsys_Project_mm_interconnect_10
		port map (
			clk_100_clk_clk                                              => m2_ddr2_memory_afi_half_clk_clk,                                            --                                            clk_100_clk.clk
			COMM_Pedreiro_v1_01_F_reset_sink_reset_bridge_in_reset_reset => rst_controller_007_reset_out_reset,                                         -- COMM_Pedreiro_v1_01_F_reset_sink_reset_bridge_in_reset.reset
			dma_comm_6_left_reset_n_reset_bridge_in_reset_reset          => rst_controller_008_reset_out_reset,                                         --          dma_comm_6_left_reset_n_reset_bridge_in_reset.reset
			dma_comm_6_left_mm_write_address                             => dma_comm_6_left_mm_write_address,                                           --                               dma_comm_6_left_mm_write.address
			dma_comm_6_left_mm_write_waitrequest                         => dma_comm_6_left_mm_write_waitrequest,                                       --                                                       .waitrequest
			dma_comm_6_left_mm_write_byteenable                          => dma_comm_6_left_mm_write_byteenable,                                        --                                                       .byteenable
			dma_comm_6_left_mm_write_write                               => dma_comm_6_left_mm_write_write,                                             --                                                       .write
			dma_comm_6_left_mm_write_writedata                           => dma_comm_6_left_mm_write_writedata,                                         --                                                       .writedata
			COMM_Pedreiro_v1_01_F_avalon_slave_L_buffer_address          => mm_interconnect_10_comm_pedreiro_v1_01_f_avalon_slave_l_buffer_address,     --            COMM_Pedreiro_v1_01_F_avalon_slave_L_buffer.address
			COMM_Pedreiro_v1_01_F_avalon_slave_L_buffer_write            => mm_interconnect_10_comm_pedreiro_v1_01_f_avalon_slave_l_buffer_write,       --                                                       .write
			COMM_Pedreiro_v1_01_F_avalon_slave_L_buffer_writedata        => mm_interconnect_10_comm_pedreiro_v1_01_f_avalon_slave_l_buffer_writedata,   --                                                       .writedata
			COMM_Pedreiro_v1_01_F_avalon_slave_L_buffer_waitrequest      => mm_interconnect_10_comm_pedreiro_v1_01_f_avalon_slave_l_buffer_waitrequest  --                                                       .waitrequest
		);

	mm_interconnect_11 : component MebX_Qsys_Project_mm_interconnect_11
		port map (
			clk_100_clk_clk                                              => m2_ddr2_memory_afi_half_clk_clk,                                            --                                            clk_100_clk.clk
			COMM_Pedreiro_v1_01_A_reset_sink_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                                         -- COMM_Pedreiro_v1_01_A_reset_sink_reset_bridge_in_reset.reset
			dma_comm_1_right_reset_n_reset_bridge_in_reset_reset         => rst_controller_008_reset_out_reset,                                         --         dma_comm_1_right_reset_n_reset_bridge_in_reset.reset
			dma_comm_1_right_mm_write_address                            => dma_comm_1_right_mm_write_address,                                          --                              dma_comm_1_right_mm_write.address
			dma_comm_1_right_mm_write_waitrequest                        => dma_comm_1_right_mm_write_waitrequest,                                      --                                                       .waitrequest
			dma_comm_1_right_mm_write_byteenable                         => dma_comm_1_right_mm_write_byteenable,                                       --                                                       .byteenable
			dma_comm_1_right_mm_write_write                              => dma_comm_1_right_mm_write_write,                                            --                                                       .write
			dma_comm_1_right_mm_write_writedata                          => dma_comm_1_right_mm_write_writedata,                                        --                                                       .writedata
			COMM_Pedreiro_v1_01_A_avalon_slave_R_buffer_address          => mm_interconnect_11_comm_pedreiro_v1_01_a_avalon_slave_r_buffer_address,     --            COMM_Pedreiro_v1_01_A_avalon_slave_R_buffer.address
			COMM_Pedreiro_v1_01_A_avalon_slave_R_buffer_write            => mm_interconnect_11_comm_pedreiro_v1_01_a_avalon_slave_r_buffer_write,       --                                                       .write
			COMM_Pedreiro_v1_01_A_avalon_slave_R_buffer_writedata        => mm_interconnect_11_comm_pedreiro_v1_01_a_avalon_slave_r_buffer_writedata,   --                                                       .writedata
			COMM_Pedreiro_v1_01_A_avalon_slave_R_buffer_waitrequest      => mm_interconnect_11_comm_pedreiro_v1_01_a_avalon_slave_r_buffer_waitrequest  --                                                       .waitrequest
		);

	mm_interconnect_12 : component MebX_Qsys_Project_mm_interconnect_12
		port map (
			clk_100_clk_clk                                              => m2_ddr2_memory_afi_half_clk_clk,                                            --                                            clk_100_clk.clk
			COMM_Pedreiro_v1_01_B_reset_sink_reset_bridge_in_reset_reset => rst_controller_003_reset_out_reset,                                         -- COMM_Pedreiro_v1_01_B_reset_sink_reset_bridge_in_reset.reset
			dma_comm_2_right_reset_n_reset_bridge_in_reset_reset         => rst_controller_008_reset_out_reset,                                         --         dma_comm_2_right_reset_n_reset_bridge_in_reset.reset
			dma_comm_2_right_mm_write_address                            => dma_comm_2_right_mm_write_address,                                          --                              dma_comm_2_right_mm_write.address
			dma_comm_2_right_mm_write_waitrequest                        => dma_comm_2_right_mm_write_waitrequest,                                      --                                                       .waitrequest
			dma_comm_2_right_mm_write_byteenable                         => dma_comm_2_right_mm_write_byteenable,                                       --                                                       .byteenable
			dma_comm_2_right_mm_write_write                              => dma_comm_2_right_mm_write_write,                                            --                                                       .write
			dma_comm_2_right_mm_write_writedata                          => dma_comm_2_right_mm_write_writedata,                                        --                                                       .writedata
			COMM_Pedreiro_v1_01_B_avalon_slave_R_buffer_address          => mm_interconnect_12_comm_pedreiro_v1_01_b_avalon_slave_r_buffer_address,     --            COMM_Pedreiro_v1_01_B_avalon_slave_R_buffer.address
			COMM_Pedreiro_v1_01_B_avalon_slave_R_buffer_write            => mm_interconnect_12_comm_pedreiro_v1_01_b_avalon_slave_r_buffer_write,       --                                                       .write
			COMM_Pedreiro_v1_01_B_avalon_slave_R_buffer_writedata        => mm_interconnect_12_comm_pedreiro_v1_01_b_avalon_slave_r_buffer_writedata,   --                                                       .writedata
			COMM_Pedreiro_v1_01_B_avalon_slave_R_buffer_waitrequest      => mm_interconnect_12_comm_pedreiro_v1_01_b_avalon_slave_r_buffer_waitrequest  --                                                       .waitrequest
		);

	mm_interconnect_13 : component MebX_Qsys_Project_mm_interconnect_13
		port map (
			clk_100_clk_clk                                              => m2_ddr2_memory_afi_half_clk_clk,                                            --                                            clk_100_clk.clk
			COMM_Pedreiro_v1_01_C_reset_sink_reset_bridge_in_reset_reset => rst_controller_004_reset_out_reset,                                         -- COMM_Pedreiro_v1_01_C_reset_sink_reset_bridge_in_reset.reset
			dma_comm_3_right_reset_n_reset_bridge_in_reset_reset         => rst_controller_008_reset_out_reset,                                         --         dma_comm_3_right_reset_n_reset_bridge_in_reset.reset
			dma_comm_3_right_mm_write_address                            => dma_comm_3_right_mm_write_address,                                          --                              dma_comm_3_right_mm_write.address
			dma_comm_3_right_mm_write_waitrequest                        => dma_comm_3_right_mm_write_waitrequest,                                      --                                                       .waitrequest
			dma_comm_3_right_mm_write_byteenable                         => dma_comm_3_right_mm_write_byteenable,                                       --                                                       .byteenable
			dma_comm_3_right_mm_write_write                              => dma_comm_3_right_mm_write_write,                                            --                                                       .write
			dma_comm_3_right_mm_write_writedata                          => dma_comm_3_right_mm_write_writedata,                                        --                                                       .writedata
			COMM_Pedreiro_v1_01_C_avalon_slave_R_buffer_address          => mm_interconnect_13_comm_pedreiro_v1_01_c_avalon_slave_r_buffer_address,     --            COMM_Pedreiro_v1_01_C_avalon_slave_R_buffer.address
			COMM_Pedreiro_v1_01_C_avalon_slave_R_buffer_write            => mm_interconnect_13_comm_pedreiro_v1_01_c_avalon_slave_r_buffer_write,       --                                                       .write
			COMM_Pedreiro_v1_01_C_avalon_slave_R_buffer_writedata        => mm_interconnect_13_comm_pedreiro_v1_01_c_avalon_slave_r_buffer_writedata,   --                                                       .writedata
			COMM_Pedreiro_v1_01_C_avalon_slave_R_buffer_waitrequest      => mm_interconnect_13_comm_pedreiro_v1_01_c_avalon_slave_r_buffer_waitrequest  --                                                       .waitrequest
		);

	mm_interconnect_14 : component MebX_Qsys_Project_mm_interconnect_14
		port map (
			clk_100_clk_clk                                              => m2_ddr2_memory_afi_half_clk_clk,                                            --                                            clk_100_clk.clk
			COMM_Pedreiro_v1_01_D_reset_sink_reset_bridge_in_reset_reset => rst_controller_005_reset_out_reset,                                         -- COMM_Pedreiro_v1_01_D_reset_sink_reset_bridge_in_reset.reset
			dma_comm_4_right_reset_n_reset_bridge_in_reset_reset         => rst_controller_008_reset_out_reset,                                         --         dma_comm_4_right_reset_n_reset_bridge_in_reset.reset
			dma_comm_4_right_mm_write_address                            => dma_comm_4_right_mm_write_address,                                          --                              dma_comm_4_right_mm_write.address
			dma_comm_4_right_mm_write_waitrequest                        => dma_comm_4_right_mm_write_waitrequest,                                      --                                                       .waitrequest
			dma_comm_4_right_mm_write_byteenable                         => dma_comm_4_right_mm_write_byteenable,                                       --                                                       .byteenable
			dma_comm_4_right_mm_write_write                              => dma_comm_4_right_mm_write_write,                                            --                                                       .write
			dma_comm_4_right_mm_write_writedata                          => dma_comm_4_right_mm_write_writedata,                                        --                                                       .writedata
			COMM_Pedreiro_v1_01_D_avalon_slave_R_buffer_address          => mm_interconnect_14_comm_pedreiro_v1_01_d_avalon_slave_r_buffer_address,     --            COMM_Pedreiro_v1_01_D_avalon_slave_R_buffer.address
			COMM_Pedreiro_v1_01_D_avalon_slave_R_buffer_write            => mm_interconnect_14_comm_pedreiro_v1_01_d_avalon_slave_r_buffer_write,       --                                                       .write
			COMM_Pedreiro_v1_01_D_avalon_slave_R_buffer_writedata        => mm_interconnect_14_comm_pedreiro_v1_01_d_avalon_slave_r_buffer_writedata,   --                                                       .writedata
			COMM_Pedreiro_v1_01_D_avalon_slave_R_buffer_waitrequest      => mm_interconnect_14_comm_pedreiro_v1_01_d_avalon_slave_r_buffer_waitrequest  --                                                       .waitrequest
		);

	mm_interconnect_15 : component MebX_Qsys_Project_mm_interconnect_15
		port map (
			clk_100_clk_clk                                              => m2_ddr2_memory_afi_half_clk_clk,                                            --                                            clk_100_clk.clk
			COMM_Pedreiro_v1_01_E_reset_sink_reset_bridge_in_reset_reset => rst_controller_006_reset_out_reset,                                         -- COMM_Pedreiro_v1_01_E_reset_sink_reset_bridge_in_reset.reset
			dma_comm_5_right_reset_n_reset_bridge_in_reset_reset         => rst_controller_008_reset_out_reset,                                         --         dma_comm_5_right_reset_n_reset_bridge_in_reset.reset
			dma_comm_5_right_mm_write_address                            => dma_comm_5_right_mm_write_address,                                          --                              dma_comm_5_right_mm_write.address
			dma_comm_5_right_mm_write_waitrequest                        => dma_comm_5_right_mm_write_waitrequest,                                      --                                                       .waitrequest
			dma_comm_5_right_mm_write_byteenable                         => dma_comm_5_right_mm_write_byteenable,                                       --                                                       .byteenable
			dma_comm_5_right_mm_write_write                              => dma_comm_5_right_mm_write_write,                                            --                                                       .write
			dma_comm_5_right_mm_write_writedata                          => dma_comm_5_right_mm_write_writedata,                                        --                                                       .writedata
			COMM_Pedreiro_v1_01_E_avalon_slave_R_buffer_address          => mm_interconnect_15_comm_pedreiro_v1_01_e_avalon_slave_r_buffer_address,     --            COMM_Pedreiro_v1_01_E_avalon_slave_R_buffer.address
			COMM_Pedreiro_v1_01_E_avalon_slave_R_buffer_write            => mm_interconnect_15_comm_pedreiro_v1_01_e_avalon_slave_r_buffer_write,       --                                                       .write
			COMM_Pedreiro_v1_01_E_avalon_slave_R_buffer_writedata        => mm_interconnect_15_comm_pedreiro_v1_01_e_avalon_slave_r_buffer_writedata,   --                                                       .writedata
			COMM_Pedreiro_v1_01_E_avalon_slave_R_buffer_waitrequest      => mm_interconnect_15_comm_pedreiro_v1_01_e_avalon_slave_r_buffer_waitrequest  --                                                       .waitrequest
		);

	mm_interconnect_16 : component MebX_Qsys_Project_mm_interconnect_16
		port map (
			clk_100_clk_clk                                              => m2_ddr2_memory_afi_half_clk_clk,                                            --                                            clk_100_clk.clk
			COMM_Pedreiro_v1_01_F_reset_sink_reset_bridge_in_reset_reset => rst_controller_007_reset_out_reset,                                         -- COMM_Pedreiro_v1_01_F_reset_sink_reset_bridge_in_reset.reset
			dma_comm_6_right_reset_n_reset_bridge_in_reset_reset         => rst_controller_008_reset_out_reset,                                         --         dma_comm_6_right_reset_n_reset_bridge_in_reset.reset
			dma_comm_6_right_mm_write_address                            => dma_comm_6_right_mm_write_address,                                          --                              dma_comm_6_right_mm_write.address
			dma_comm_6_right_mm_write_waitrequest                        => dma_comm_6_right_mm_write_waitrequest,                                      --                                                       .waitrequest
			dma_comm_6_right_mm_write_byteenable                         => dma_comm_6_right_mm_write_byteenable,                                       --                                                       .byteenable
			dma_comm_6_right_mm_write_write                              => dma_comm_6_right_mm_write_write,                                            --                                                       .write
			dma_comm_6_right_mm_write_writedata                          => dma_comm_6_right_mm_write_writedata,                                        --                                                       .writedata
			COMM_Pedreiro_v1_01_F_avalon_slave_R_buffer_address          => mm_interconnect_16_comm_pedreiro_v1_01_f_avalon_slave_r_buffer_address,     --            COMM_Pedreiro_v1_01_F_avalon_slave_R_buffer.address
			COMM_Pedreiro_v1_01_F_avalon_slave_R_buffer_write            => mm_interconnect_16_comm_pedreiro_v1_01_f_avalon_slave_r_buffer_write,       --                                                       .write
			COMM_Pedreiro_v1_01_F_avalon_slave_R_buffer_writedata        => mm_interconnect_16_comm_pedreiro_v1_01_f_avalon_slave_r_buffer_writedata,   --                                                       .writedata
			COMM_Pedreiro_v1_01_F_avalon_slave_R_buffer_waitrequest      => mm_interconnect_16_comm_pedreiro_v1_01_f_avalon_slave_r_buffer_waitrequest  --                                                       .waitrequest
		);

	irq_mapper : component MebX_Qsys_Project_irq_mapper
		port map (
			clk            => m2_ddr2_memory_afi_half_clk_clk,    --        clk.clk
			reset          => rst_controller_012_reset_out_reset, --  clk_reset.reset
			receiver0_irq  => irq_mapper_receiver0_irq,           --  receiver0.irq
			receiver1_irq  => irq_mapper_receiver1_irq,           --  receiver1.irq
			receiver2_irq  => irq_mapper_receiver2_irq,           --  receiver2.irq
			receiver3_irq  => irq_mapper_receiver3_irq,           --  receiver3.irq
			receiver4_irq  => irq_mapper_receiver4_irq,           --  receiver4.irq
			receiver5_irq  => irq_mapper_receiver5_irq,           --  receiver5.irq
			receiver6_irq  => irq_mapper_receiver6_irq,           --  receiver6.irq
			receiver7_irq  => irq_mapper_receiver7_irq,           --  receiver7.irq
			receiver8_irq  => irq_mapper_receiver8_irq,           --  receiver8.irq
			receiver9_irq  => irq_mapper_receiver9_irq,           --  receiver9.irq
			receiver10_irq => irq_mapper_receiver10_irq,          -- receiver10.irq
			receiver11_irq => irq_mapper_receiver11_irq,          -- receiver11.irq
			receiver12_irq => irq_mapper_receiver12_irq,          -- receiver12.irq
			receiver13_irq => irq_mapper_receiver13_irq,          -- receiver13.irq
			receiver14_irq => irq_mapper_receiver14_irq,          -- receiver14.irq
			receiver15_irq => irq_mapper_receiver15_irq,          -- receiver15.irq
			receiver16_irq => irq_mapper_receiver16_irq,          -- receiver16.irq
			receiver17_irq => irq_mapper_receiver17_irq,          -- receiver17.irq
			receiver18_irq => irq_mapper_receiver18_irq,          -- receiver18.irq
			receiver19_irq => irq_mapper_receiver19_irq,          -- receiver19.irq
			receiver20_irq => irq_mapper_receiver20_irq,          -- receiver20.irq
			receiver21_irq => irq_mapper_receiver21_irq,          -- receiver21.irq
			receiver22_irq => irq_mapper_receiver22_irq,          -- receiver22.irq
			receiver23_irq => irq_mapper_receiver23_irq,          -- receiver23.irq
			receiver24_irq => irq_mapper_receiver24_irq,          -- receiver24.irq
			receiver25_irq => irq_mapper_receiver25_irq,          -- receiver25.irq
			receiver26_irq => irq_mapper_receiver26_irq,          -- receiver26.irq
			receiver27_irq => irq_mapper_receiver27_irq,          -- receiver27.irq
			receiver28_irq => irq_mapper_receiver28_irq,          -- receiver28.irq
			receiver29_irq => irq_mapper_receiver29_irq,          -- receiver29.irq
			receiver30_irq => irq_mapper_receiver30_irq,          -- receiver30.irq
			receiver31_irq => irq_mapper_receiver31_irq,          -- receiver31.irq
			sender_irq     => nios2_gen2_0_irq_irq                --     sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk50_clk,                          --       receiver_clk.clk
			sender_clk     => m2_ddr2_memory_afi_half_clk_clk,    --         sender_clk.clk
			receiver_reset => rst_controller_009_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_012_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver21_irq           --             sender.irq
		);

	irq_synchronizer_001 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk50_clk,                          --       receiver_clk.clk
			sender_clk     => m2_ddr2_memory_afi_half_clk_clk,    --         sender_clk.clk
			receiver_reset => rst_controller_009_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_012_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_001_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver22_irq           --             sender.irq
		);

	irq_synchronizer_002 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk50_clk,                          --       receiver_clk.clk
			sender_clk     => m2_ddr2_memory_afi_half_clk_clk,    --         sender_clk.clk
			receiver_reset => rst_controller_013_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_012_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_002_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver23_irq           --             sender.irq
		);

	irq_synchronizer_003 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk50_clk,                          --       receiver_clk.clk
			sender_clk     => m2_ddr2_memory_afi_half_clk_clk,    --         sender_clk.clk
			receiver_reset => rst_controller_014_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_012_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_003_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver24_irq           --             sender.irq
		);

	irq_synchronizer_004 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => clk50_clk,                          --       receiver_clk.clk
			sender_clk     => m2_ddr2_memory_afi_half_clk_clk,    --         sender_clk.clk
			receiver_reset => rst_controller_014_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_012_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_004_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver31_irq           --             sender.irq
		);

	rst_controller_001 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                     -- reset_in0.reset
			reset_in1      => rst_controller_reset_source_sd_card_reset, -- reset_in1.reset
			clk            => clk50_clk,                                 --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,        -- reset_out.reset
			reset_req      => open,                                      -- (terminated)
			reset_req_in0  => '0',                                       -- (terminated)
			reset_req_in1  => '0',                                       -- (terminated)
			reset_in2      => '0',                                       -- (terminated)
			reset_req_in2  => '0',                                       -- (terminated)
			reset_in3      => '0',                                       -- (terminated)
			reset_req_in3  => '0',                                       -- (terminated)
			reset_in4      => '0',                                       -- (terminated)
			reset_req_in4  => '0',                                       -- (terminated)
			reset_in5      => '0',                                       -- (terminated)
			reset_req_in5  => '0',                                       -- (terminated)
			reset_in6      => '0',                                       -- (terminated)
			reset_req_in6  => '0',                                       -- (terminated)
			reset_in7      => '0',                                       -- (terminated)
			reset_req_in7  => '0',                                       -- (terminated)
			reset_in8      => '0',                                       -- (terminated)
			reset_req_in8  => '0',                                       -- (terminated)
			reset_in9      => '0',                                       -- (terminated)
			reset_req_in9  => '0',                                       -- (terminated)
			reset_in10     => '0',                                       -- (terminated)
			reset_req_in10 => '0',                                       -- (terminated)
			reset_in11     => '0',                                       -- (terminated)
			reset_req_in11 => '0',                                       -- (terminated)
			reset_in12     => '0',                                       -- (terminated)
			reset_req_in12 => '0',                                       -- (terminated)
			reset_in13     => '0',                                       -- (terminated)
			reset_req_in13 => '0',                                       -- (terminated)
			reset_in14     => '0',                                       -- (terminated)
			reset_req_in14 => '0',                                       -- (terminated)
			reset_in15     => '0',                                       -- (terminated)
			reset_req_in15 => '0'                                        -- (terminated)
		);

	rst_controller_002 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                      -- reset_in0.reset
			reset_in1      => rst_controller_reset_source_comm_ch1_reset, -- reset_in1.reset
			clk            => m2_ddr2_memory_afi_half_clk_clk,            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,         -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	rst_controller_003 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                      -- reset_in0.reset
			reset_in1      => rst_controller_reset_source_comm_ch2_reset, -- reset_in1.reset
			clk            => m2_ddr2_memory_afi_half_clk_clk,            --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset,         -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	rst_controller_004 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                      -- reset_in0.reset
			reset_in1      => rst_controller_reset_source_comm_ch3_reset, -- reset_in1.reset
			clk            => m2_ddr2_memory_afi_half_clk_clk,            --       clk.clk
			reset_out      => rst_controller_004_reset_out_reset,         -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	rst_controller_005 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                      -- reset_in0.reset
			reset_in1      => rst_controller_reset_source_comm_ch4_reset, -- reset_in1.reset
			clk            => m2_ddr2_memory_afi_half_clk_clk,            --       clk.clk
			reset_out      => rst_controller_005_reset_out_reset,         -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	rst_controller_006 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                      -- reset_in0.reset
			reset_in1      => rst_controller_reset_source_comm_ch5_reset, -- reset_in1.reset
			clk            => m2_ddr2_memory_afi_half_clk_clk,            --       clk.clk
			reset_out      => rst_controller_006_reset_out_reset,         -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	rst_controller_007 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                      -- reset_in0.reset
			reset_in1      => rst_controller_reset_source_comm_ch6_reset, -- reset_in1.reset
			clk            => m2_ddr2_memory_afi_half_clk_clk,            --       clk.clk
			reset_out      => rst_controller_007_reset_out_reset,         -- reset_out.reset
			reset_req      => open,                                       -- (terminated)
			reset_req_in0  => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	rst_controller_008 : component mebx_qsys_project_rst_controller_008
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                  -- reset_in0.reset
			clk            => m2_ddr2_memory_afi_half_clk_clk,        --       clk.clk
			reset_out      => rst_controller_008_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_008_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_009 : component mebx_qsys_project_rst_controller_009
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
			clk            => clk50_clk,                          --       clk.clk
			reset_out      => rst_controller_009_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_010 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
			reset_in1      => rst_reset_n_ports_inv,              -- reset_in1.reset
			clk            => m2_ddr2_memory_afi_half_clk_clk,    --       clk.clk
			reset_out      => rst_controller_010_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_011 : component mebx_qsys_project_rst_controller_009
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
			clk            => m1_ddr2_memory_afi_half_clk_clk,    --       clk.clk
			reset_out      => rst_controller_011_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_012 : component mebx_qsys_project_rst_controller_008
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                  -- reset_in0.reset
			clk            => m2_ddr2_memory_afi_half_clk_clk,        --       clk.clk
			reset_out      => rst_controller_012_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_012_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_013 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                   -- reset_in0.reset
			reset_in1      => rst_controller_reset_source_rs232_reset, -- reset_in1.reset
			clk            => clk50_clk,                               --       clk.clk
			reset_out      => rst_controller_013_reset_out_reset,      -- reset_out.reset
			reset_req      => open,                                    -- (terminated)
			reset_req_in0  => '0',                                     -- (terminated)
			reset_req_in1  => '0',                                     -- (terminated)
			reset_in2      => '0',                                     -- (terminated)
			reset_req_in2  => '0',                                     -- (terminated)
			reset_in3      => '0',                                     -- (terminated)
			reset_req_in3  => '0',                                     -- (terminated)
			reset_in4      => '0',                                     -- (terminated)
			reset_req_in4  => '0',                                     -- (terminated)
			reset_in5      => '0',                                     -- (terminated)
			reset_req_in5  => '0',                                     -- (terminated)
			reset_in6      => '0',                                     -- (terminated)
			reset_req_in6  => '0',                                     -- (terminated)
			reset_in7      => '0',                                     -- (terminated)
			reset_req_in7  => '0',                                     -- (terminated)
			reset_in8      => '0',                                     -- (terminated)
			reset_req_in8  => '0',                                     -- (terminated)
			reset_in9      => '0',                                     -- (terminated)
			reset_req_in9  => '0',                                     -- (terminated)
			reset_in10     => '0',                                     -- (terminated)
			reset_req_in10 => '0',                                     -- (terminated)
			reset_in11     => '0',                                     -- (terminated)
			reset_req_in11 => '0',                                     -- (terminated)
			reset_in12     => '0',                                     -- (terminated)
			reset_req_in12 => '0',                                     -- (terminated)
			reset_in13     => '0',                                     -- (terminated)
			reset_req_in13 => '0',                                     -- (terminated)
			reset_in14     => '0',                                     -- (terminated)
			reset_req_in14 => '0',                                     -- (terminated)
			reset_in15     => '0',                                     -- (terminated)
			reset_req_in15 => '0'                                      -- (terminated)
		);

	rst_controller_014 : component mebx_qsys_project_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,                  -- reset_in0.reset
			reset_in1      => rst_controller_reset_source_sync_reset, -- reset_in1.reset
			clk            => clk50_clk,                              --       clk.clk
			reset_out      => rst_controller_014_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_015 : component mebx_qsys_project_rst_controller_009
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
			clk            => m2_ddr2_memory_afi_clk_clk,         --       clk.clk
			reset_out      => rst_controller_015_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_016 : component mebx_qsys_project_rst_controller_009
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rst_reset_n_ports_inv,              -- reset_in0.reset
			clk            => m1_ddr2_memory_afi_clk_clk,         --       clk.clk
			reset_out      => rst_controller_016_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_reset_n_ports_inv <= not rst_reset_n;

	mm_interconnect_0_m2_ddr2_memory_avl_inv <= not m2_ddr2_memory_avl_waitrequest;

	mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_2_m1_ddr2_i2c_sda_s1_write_ports_inv <= not mm_interconnect_2_m1_ddr2_i2c_sda_s1_write;

	mm_interconnect_2_m1_ddr2_i2c_scl_s1_write_ports_inv <= not mm_interconnect_2_m1_ddr2_i2c_scl_s1_write;

	mm_interconnect_2_pio_led_s1_write_ports_inv <= not mm_interconnect_2_pio_led_s1_write;

	mm_interconnect_2_timer_1ms_s1_write_ports_inv <= not mm_interconnect_2_timer_1ms_s1_write;

	mm_interconnect_2_timer_1us_s1_write_ports_inv <= not mm_interconnect_2_timer_1us_s1_write;

	mm_interconnect_2_temp_scl_s1_write_ports_inv <= not mm_interconnect_2_temp_scl_s1_write;

	mm_interconnect_2_temp_sda_s1_write_ports_inv <= not mm_interconnect_2_temp_sda_s1_write;

	mm_interconnect_2_m2_ddr2_i2c_sda_s1_write_ports_inv <= not mm_interconnect_2_m2_ddr2_i2c_sda_s1_write;

	mm_interconnect_2_m2_ddr2_i2c_scl_s1_write_ports_inv <= not mm_interconnect_2_m2_ddr2_i2c_scl_s1_write;

	mm_interconnect_2_csense_sdi_s1_write_ports_inv <= not mm_interconnect_2_csense_sdi_s1_write;

	mm_interconnect_2_csense_sck_s1_write_ports_inv <= not mm_interconnect_2_csense_sck_s1_write;

	mm_interconnect_2_csense_cs_n_s1_write_ports_inv <= not mm_interconnect_2_csense_cs_n_s1_write;

	mm_interconnect_2_csense_adc_fo_s1_write_ports_inv <= not mm_interconnect_2_csense_adc_fo_s1_write;

	mm_interconnect_2_pio_led_painel_s1_write_ports_inv <= not mm_interconnect_2_pio_led_painel_s1_write;

	mm_interconnect_2_rtcc_sdi_s1_write_ports_inv <= not mm_interconnect_2_rtcc_sdi_s1_write;

	mm_interconnect_2_rtcc_sck_s1_write_ports_inv <= not mm_interconnect_2_rtcc_sck_s1_write;

	mm_interconnect_2_rtcc_cs_n_s1_write_ports_inv <= not mm_interconnect_2_rtcc_cs_n_s1_write;

	mm_interconnect_2_rs232_uart_s1_read_ports_inv <= not mm_interconnect_2_rs232_uart_s1_read;

	mm_interconnect_2_rs232_uart_s1_write_ports_inv <= not mm_interconnect_2_rs232_uart_s1_write;

	mm_interconnect_2_pio_ctrl_io_lvds_s1_write_ports_inv <= not mm_interconnect_2_pio_ctrl_io_lvds_s1_write;

	mm_interconnect_3_m1_ddr2_memory_avl_inv <= not m1_ddr2_memory_avl_waitrequest;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_008_reset_out_reset_ports_inv <= not rst_controller_008_reset_out_reset;

	rst_controller_009_reset_out_reset_ports_inv <= not rst_controller_009_reset_out_reset;

	rst_controller_012_reset_out_reset_ports_inv <= not rst_controller_012_reset_out_reset;

	rst_controller_013_reset_out_reset_ports_inv <= not rst_controller_013_reset_out_reset;

end architecture rtl; -- of MebX_Qsys_Project
