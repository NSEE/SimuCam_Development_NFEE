// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
JX8xeTO4VIu71/t3q1YzOjz8IJa1w3pWjtnOQvHFIUQe0qX15ja+dSqVX/qZAlcJgY/CZ1BVR7kh
keOD+Hct2g61UWtbqTfkE61/UIrgbLAQU4V+xkL6ZGkXVgfWt48OkwbEGVdBrbzPoJDbdX6+zkJf
K5PHVUfWZg7cOHuW2+KxS5RnUih2S+LtJahmjkhXm7GraoPEAGuGsRNCC/2ME/ZOobW5ZO+kyh7a
0erV76E0VKcuIB1I1dz4ldfqFY277Dsx/60Zo9p3+lO7vOcABIfoEcSusVFTVZUFmzG4ZhSR6MCR
3+mn2OUl/1a/ueb3c9e2FNsTo9we59AtnZpzWQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5616)
yCLeYYtxHKOSnP+qktFIV3ymsPW1vG7IIl7kCwN+IW4nYt+sItC16KwR6F73w8cGF7SBmALEhMj4
T0uQiyIYSylTxLbrpa2MNAddFaKMMDmWTUzmB9v4uX0Jl3KH3wfBo8Y6R5aqEPmR6GJItORmZzrp
ozC4qU++YTqezJwOyjVzeWVsORiZ2uZg3q8P+NHt/AtR4cNmVtA1PIqzC3Hq7xYPs++FehvcJAJ8
ltbddk7Wwe/aGE1H19YQAmLriYWGwdVjsCqCKzobUk7hUZHeB/DDuyte1a2eyL5yWBUUFeElxdZT
Umyq4W4IRaIhEjHI/3qEASLyc4vV1uIqMqE1qxpK+f+2vyCQtKl9BqpXG2CyBBXm1KreW3uarbkX
rUf0BrqFUPF9+RdlQU4hsJQYvJRyML5IDd4Gv36Hfw852t9l1prMZxg8PrBtIJ5UJjFgd/xrix98
KECT4qkeIBv3D33ZngkFfdms9y+R/u7zAsfY0flqPDy1oEA56XCQClJQK8z8sYSzmkGttBSWDSs5
fe4z7ol7fg7S9wU1lP7ExngRrY/BbI+AXPtQEMJMz2qqU6QJ55sjZ38pw3gDk6hulGcjE7Y0IGDe
lAp17J/Qoe1S+O+jvSHc1BjdvCsFRWQjJDDOSdyE9LDojUp+saskE5uKLQG6gaWwzWrrlljk+s/z
91xeUtWPa9M7sBOhk11c9QjijjrR+lzsfrv7L/hqesIhHyl1FI4W2P20lHRMwBznP8acRhR0JTIT
jKw1X+1aS/Rnn38VYst1Ogc0OlRncT38m9w/dEjoTV4L59/iCUGltC1PViv2BHmIee2U+NGmGGew
fTjcS/MnZzsZ5WO0+GZYexwnV4fCLFPL/z+bJbOAgPJdcVMpFTSz7Hu82q3zyOJEb4OSh07kALCG
di8xLAo072JWRK6XBudHAwgHTOmkeRuqcD+qB0TcXxzWDFvN9baMkZgp0NgQmvYhrHaMNsmXUY7C
AsSAsS8pIQxZHRsi423VHYIUsYE5Bin3m6TUztmbTMn50Q1a0E9JEnYIoXaaOQJB0RY0Laythab7
xKey5OL+bUignhu9/d4FORLpygccmd4rrTKORj0WE12XF3nX4ZINEGYEWsvuysEJj9bLVwYuq+9n
bevGGmnuc/IogsP/N8sVGUvcT/N5pnCPkgHzT2IM1qmRd13H8yBRSX9W1ljQeUDbkqoyrUTAePfl
xO2TJM3JHhPJhmm1ZMJyJBHF7oMuFNo9wawq/jP4vjmFOu+5Ids6/JxjkLXb2ZEUzrnwQxoY8mIn
g9iXuZBUwXC8073AZMwutL4mnDUppCONu2Nqji+Rs2AJ6pU/KkRXusvOiifVrCotXvL9T9BBi8X1
MxWhE66NeSqTPAJtKIHKjQQV4ubyI1mIc77BlStza2pQ+UZpk9PQ9rdQO4+8GEV6MFFTPTyOzD+e
lLVP27PUhpJMKakfivtn6zDbUy414Jfjnzr341FpKcf/6voNALssqFBsCuhSVuexfVYEuNYLf1Cu
P3c3+y8YZU3rdzbReec6uJkzMchH8HggM+7ihf0LQ9qNL8XMcIjuR0QMlDS7IJa9YClBKddvg4e+
puztONslsTPXMLRjE7JmPUTUKcEDYI9ratnig+qmbZ/eNic3Q1NnZglXXcSNnEyrQiQWg4l3KPof
S7jXOUPOz2A82pyR5VnWbh0UuZgPM2Pbm5OmfhNioKWrtMttbtMrJYn/ew35bKx5evea4SG87MHp
LHlvD1VtlbOrPzhneBlVt83xbLpenhviRWO01MhOeZqyhCSPl5nvoPLbwDi+I8/AXJCZvKivs6ab
X3zNJy6oohdeJVr186aG5rnpHsNoo2iLPivjuSRTQth7G3jTnGkdgIo5DzxC2gMU1uixDsSxuchI
6GRU6ero89Eoggujv80uwyyv45vTlaRYv1ep4mblRfeUIdjdr/gQCMy8fdlxJ8jjDNvr4my3SU33
TxTcW5Ck6MiXfRBx2b4Xu3xycgF8e2u71zImNxK4TrvPp5qAmXMTb46bJxb33+yscNbohwbk5p2B
dJLVrOKEmAIoZzUfGXIvgoPpkQQ8pd0rvOkrYs3nx5oqeQ6ppLd6NF4Tc0+FGoJc0Em99MHSB3QQ
SPLlfXybleRo+fE3UhIn4ztzEfZEF7cF2+L27pRaNEFVcV8aDil03ciiR06aFJZts5k4kB+4RVjk
yVOQUHFz0URisoNUX8rzC/+jKSJ4cgkxErlRBVvWp29DdBmZ+U5Cdztaao211m/tAEEBCA5MnYO6
GWl34KNZ3MWrK4CBJnzcN1+tQzUtlunVKuwD3h6ZbHDPPt+SsSKyP46mqDD+ZLS4lyE8u96jojgq
rJkNzCxrzuazqYrtWDKw5pr5rmtab44O1ZQ4XojArQaiAPY3KA4jO3tU+gNy94dHUPPdbMwXWW6G
h8XPjZHabGNW/YL1Cjo+v4QbbHgRY4LkYD656cCbrVlKYRbgLAUL1dKXXNgTywHbfHHPxGQv2xy2
PBoiF6Mbrh4klq6XNdat78JvNLRz5ItY4DrCROHbw4lGyfui8mPP6JcuyoZ9U4APVitLWHM3i4Kj
CEvLXAYDtKLtr1WyRMIK0kVlp7mUVLwXedHrlGc1qmwdAHPrufvVfiNtrsOV0FJxEcZlFSQrIEZ1
0yA/wgqhVPOLgjpoSYJK12yFq0zGRynChU+Oszf+gyUma5kvXrfYM0erSq4fsxAM/uINT5wUKAVu
sbhZw39NO83sinYadW2gjgKt3WoQHIkFTCnrEq0kDyP0dkRCcgFwMmU4ArJh5YHywK7KV9Lxl3wm
Vtvp18pe8OxSoNtAtjMSRHSA/yU8DYTQq8VmUneGHPcMrdA3XkvH3Xhpv3rFNcDeNEYOhGaHcV6L
4iFUJECXQE1CvYMT+BDXCTogAXpwl6ertz/DIJEgXMUqz8GiassWN7Tem33UwkhqeeDLNMgs4bXA
uGzmrNKSRhh2lro3EuPNnPRaL95gku48AXOSbzNigZ7LpfqQxCpNGlBwDBVSVuT9Qx8Zl1nHeqJD
v+KJZWyteebJQOwT9a35VoAQcLrtV2djIJYZqpuKetfvca2s1IIFgwLeiRXEZD1SiwL2tjg/As7E
C5CX0MynsaUxFxZZIMO12ETngOKAOl9IaqgYeI2yd/wiSqg2LqXU7RhPD0wqxkgoqOiTzc/LhBN7
PvoQsQAh0h1BIW84DxAMj3gvweLqE94zf4QWipxBLzX237NkGWcRTvN+JjxMJxCyVTKe5GCW0u+j
y4+u+6pXD3flyMb2KVG1CFtmGA6OGd/yiycvLcGCJXEFOHsZma+ttS/saIUxKN5hT+6LmJkTdkVc
DnYwThC3JRnp4uD8IoMOshkAiEd2ogSOHsRqjkVBWCnS85gsBaPSw/StIwbWHXtEsVIPcaIekM69
hQW74maHqMUgtugqYPdUAuyhYtD0e4QcK41c1MXlcn8kJoBpwAF75TtG/tEe2zZxKp9WnEI4h60I
EnnQkjoEysG0Vh1neLGXH4wD41r/inEX9L0QQwOca6ZzDdT71bzD//KfR5h2GDfvnhRBlOCn9Uyp
GnkYGUh1DZfFqGNlkrOatp9gBrF6XWRjbFJ8pIrtGWZo1lA+ClW642eZjAKAhcc3QGNisBqz3tCy
tjBtse1G5+DmcMAHvaD0WxQ+6FDP4Db40HzZfFFUims8Vss2aarVBH+dc2M/2pSvkfgAegUZDcxf
CN7fX2rIkuwH6etVpZDUDKtMXOuJrGhJtoI6QzmogmiGagwDl53NoGRu+8QP1nBxxjmbQv/Y1qpj
6d+AQXtoPfJQ00A5IZmYU60ewbytUHY7OeSjIrZM2+6W9LjenPHYCHr6a/bTZIFQoaHe6dgiNoYy
6tSCHK1lFkYoUNmSFtikPao0dUDesqm02/sbjfDj+dkC1g/XXDJXRtzkR/lOh6EfJ/9QWM/bQP5D
m+Mc4zESuenCs98Frb1O0n3YN8zXNoGO0uGtr98nEgCvxPOm3Bm4pW6a2XwNcVs3bB+ivmOz/KMV
+OArdHWeOwtOqbDn/teew8vbwZj+nm6qho7Spi+aLT7ie4FrCFaTAb20tGuZcA7DMcxpR+DAMvMw
+usXJ2dtjPWftk3Tk2jPbGHVGllcap1xoyWl9z1hSffdURyunhdqv+5sy7RC38qgLj1knmz+vnv6
z+P5hkrY7tK8lx8iZ5+RT5jtcQa3IN/9vo9ioHhrjYpaSMuF1v0rokFgYfzSnywQcGFiz0z0aFpD
mZQWpoabktKTMwiR+oLo9HwGwsW6lhenVdn0qifroQZ5hwVZsY19jkQGBOulBRg75+KDfWeHai5Y
7rSc2OXkTf6NML9E3X/PLMMrLbb5QR99/rcUWU2KWL9Glh40F14Qz3+4LlC+Xk7AndXt5g3n56f3
PX0ISf7NKFyLc/eEacCCEPF6oLl23Es/GAMwcsRl++RzlQVRIUoXoyemY6M/mizP4uFDWAMolk/c
26KTvlnOJT+LrvqrbLgAEJs2T9PCqZBSOU7xtw28qJ480yZEalGycTdv0NnTe+fyp+E28AoCkXJq
hsLvfKDWVvV56xb0nbSFSFpoweMtT4QlGh7zWwtxnPzlCud/ihGtIYsu//+KFF9anli32I0GxwCn
LxhY5ZNabrrkfe/er3WykQ74Rv0zEjiTsypy4/WmK1oef7q5e04lHCIFNs8Ixt91Lb2U0RF1a/8j
jXLF1GZXJdQVBbK8JXyfX8PlSRuSXpNYIYnmov1U4p4ZcjImKogwHezKIAnP3kGX4ugDY/kTtEbp
IcEEErSITh+jmXJbiqe5NXs1QSJfAR47whX7IWejwVmq121KdQ/4xjpMfPbUX+AaTn07yXgwogM6
M+z5GaCjAn9N+oguJH7iputKrraHqdCSW6uqlO+6FCITbrAbmPMrK4GfmV9zkRLOl62zH00v8kai
yIxKKoLOh9J/Bd/WNIQDUTxF2AMHcKiAR3kUJtV53fxNblxXrbEBU0i7o8UoWJSAqF1HXu9wfH/N
fdx0mQqoG95OV5U7noASYzybrEzJ5K6QbuZ093/b6WVzncNRQLdOQFMQV8oJr3LhNn4RlawIvftg
4BHQPmYwpFo+3XPXyvAotsdp/y5YXa/Z9AeO5lNNbMSHVDFZhWlAGWuSxr3ovNwQ4FXbVmXvpZTQ
ngq91iXBnPWHt6FimV4eN3GA1mbJ80JZpRxwb9uER45Yqq1xULzVHhKde5c3mwIrn/nnviO6uDJl
g3c+jZ8uuFJg6myf3nMFv59QYde+hBBGIWlNYyWYue4KujDDWKd/stmvNQUL2Au/rHFXUtcxhwQu
1Y0uDXF23oQ8hqyG0QdYIEvKAkoLX+dQztcF0c98rrqVFsVKKJkkWJia4JE6bZnf2pCDYYb+yUmY
sy8KqNrxgPFD6z/R2SuFPvSy061ZjvARHMxRh2vIiQ9ieGNna3cGmneSlZZzYgchOOiD90WI8mqn
ugZNt21nTOt/66WA66O4ybVcT+TXeuy0a9RkCXoIaUfULM5kjrqAIwCFns3xYiyCrEG2+St9sa9G
dszdrRMmCDR6mKrVUQGwlfscTus4+XlFxE7aXhoHUPEAeB+fUdTSg19X4SU/InnH24ziTBMTQx9Z
4OjIbnndkbsjmz2/ZOB7XsN1/dveSHrmaCTpirGWnzT+ikp7TXih32NEeY8cCiV3v6oGAxU24nwd
LVedZ8I7eYNIK/SnihewdKjfNKpCO3H23pjA+O43x07xA2XLMQg4UNQT6k8gj4MsLx9D5FXn2vgj
mGpzmv3439AQdfzlUqDwwWA+OUEcL+739mxDHQgMsV6pF9wBWragbuzWlbXi2ti7ldEfZBexHxgk
hmt1G1HufS3eVtIPuh7eJunxczT3MkW+OzRL6KJ0R/z2+ojgDOiCL/wm1KWeXcR01Q7int0hRiKt
vFZdwpFHgaES9QGJfwzhgasFk3LqSlsoOL/hDRLrWEtpz/FwKWNGOgAB5+294n3gkIMtn/0d0MIu
AF7iNxIS68ITS1zfEm6J6rqUTxscKn3p1WrfrR1f8FNWkNjmqZJsnO8AAKM7enrqndjCkcbYEs8A
bfrAn0UYdGnBYHcjpf6LMXPuYhoTLXNliYZAN5UPyMFrEgDFeDg6hLg+AylWT8pPjY5uC2DVkdUA
uvXlSzF6XySVmI0JptvKTpDFvHlgkMNkzhJDKrhfYK8y0cSytozMA38sg6E3Kv6zHjbLc11je07V
rGy5ZkWcYKDezXQuKGl59I8NpUJS2wn1RjQz5FjrzApKpLpqbW+MCGrYpUa8mletv/mX6iR/6UuY
uL/MeTyXU0OOs6ScFqeJfkY7FYQ6tdncg0d9P6f+ve0bSyoM6ndWHBSCrBBy3vWwCDCXgoFDrQtd
yY2XjBjGJHjBJlmq94FZWWYevaMjqe307uqeCr8it/7F/ROlIx5Ew9mgWbsH10w3n7HaCDkY+Dcr
ZXppWcEq53Lio23J+YGDaWPqC0nqLGZiF1QhN+gFz2rB6mve1RYmDBB2UiH9dOZIYhMy9a3b5KA8
paLrgpbRECUSlQaU6jZiJJ2Ryyphd1UJxXW6fYNEwfSttAwnG6hQYBHVuzr3fH9e5v3rBY3Nk6Ao
mde/1bVi6Z22zJYH9GIgWm1kAg+jUmSrqrtkJrbP2uQxeLS31KdSaYGlZWjEnqiJVAF35lBc6jJs
7PXU44UZdWqUJOTtnJRW7KpFFX7lkpBQyH26e7gcoCoyPVXy9FWscaJ5NqHD3cimvSPKWBIxA3t8
w4mMw4ea/z3RxRkFi27Q8qt6yWHKQpjGo8ZHt/TaMLVPANgqebTdtpsl/aawT3/VmAMbPf3Zsnpt
hDt/iRF7b+/GPg78QHYhKLIlYTebgyjUFHdC9Rv9icI9noGWg3JK+4iFgpf2vJOp35+gT+rCivA9
JipXRDW5IbsP4/I1WS2uHibV6qmAVS7fJbD/AQICfNOKy4pvusVXXR1eOZ7av0JwqR7vochuxAMM
TBEWf89idlWD1rvMRcW3++tIm68zJjBEma/s0VHII8FUNwOvI/1Hs0NIi+4bCOSsz4zJDZAyQndS
a6vv9R2xw/sdTBlvqWMYOoOG07+QYiU/osbwDneP7Ksl3FZHbHUd0D72n3HkbKNL4e0yhr4hZ3wx
KgqWPok8AX18RSeQyBlkSsYOzYEMH/2Rpqyp7AY6YWyAaWiITpairG/qyIzKTQXf8CdABKeOSaHO
RyWCLUnxATbP8Cqn48XNHiDLt1vy6TzDhix5iOGjtYy30NmT2KAmmjOI1zg6yrTNZBxeL1+/AM/X
xyt70brZhwCy/klSpEC7QiUudz9p7SXVmH1d8UloGFgyZow7HN50ufbYmUPBERwS8Zw5269bcUTL
apJLxBHWjOy8uiSRpBT8htHvrcnxgy/0B9/fvjQUmQXSYKC6lXA/TaN/sm3Zjb10twQbZZar+BWf
d/B06O8PCmRk2t8Dw9BfBQWfO8CrbFjnJTWxmB3E
`pragma protect end_protected
