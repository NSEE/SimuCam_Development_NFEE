io_in_3b_inst : io_in_3b PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig
	);
