// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.



// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// $Id: //acds/rel/18.1std/ip/merlin/altera_merlin_router/altera_merlin_router.sv.terp#1 $
// $Revision: #1 $
// $Date: 2018/07/18 $
// $Author: psgswbuild $

// -------------------------------------------------------
// Merlin Router
//
// Asserts the appropriate one-hot encoded channel based on 
// either (a) the address or (b) the dest id. The DECODER_TYPE
// parameter controls this behaviour. 0 means address decoder,
// 1 means dest id decoder.
//
// In the case of (a), it also sets the destination id.
// -------------------------------------------------------

`timescale 1 ns / 1 ns

module MebX_Qsys_Project_mm_interconnect_0_router_032_default_decode
  #(
     parameter DEFAULT_CHANNEL = 0,
               DEFAULT_WR_CHANNEL = -1,
               DEFAULT_RD_CHANNEL = -1,
               DEFAULT_DESTID = 24 
   )
  (output [390 - 386 : 0] default_destination_id,
   output [32-1 : 0] default_wr_channel,
   output [32-1 : 0] default_rd_channel,
   output [32-1 : 0] default_src_channel
  );

  assign default_destination_id = 
    DEFAULT_DESTID[390 - 386 : 0];

  generate
    if (DEFAULT_CHANNEL == -1) begin : no_default_channel_assignment
      assign default_src_channel = '0;
    end
    else begin : default_channel_assignment
      assign default_src_channel = 32'b1 << DEFAULT_CHANNEL;
    end
  endgenerate

  generate
    if (DEFAULT_RD_CHANNEL == -1) begin : no_default_rw_channel_assignment
      assign default_wr_channel = '0;
      assign default_rd_channel = '0;
    end
    else begin : default_rw_channel_assignment
      assign default_wr_channel = 32'b1 << DEFAULT_WR_CHANNEL;
      assign default_rd_channel = 32'b1 << DEFAULT_RD_CHANNEL;
    end
  endgenerate

endmodule


module MebX_Qsys_Project_mm_interconnect_0_router_032
(
    // -------------------
    // Clock & Reset
    // -------------------
    input clk,
    input reset,

    // -------------------
    // Command Sink (Input)
    // -------------------
    input                       sink_valid,
    input  [404-1 : 0]    sink_data,
    input                       sink_startofpacket,
    input                       sink_endofpacket,
    output                      sink_ready,

    // -------------------
    // Command Source (Output)
    // -------------------
    output                          src_valid,
    output reg [404-1    : 0] src_data,
    output reg [32-1 : 0] src_channel,
    output                          src_startofpacket,
    output                          src_endofpacket,
    input                           src_ready
);

    // -------------------------------------------------------
    // Local parameters and variables
    // -------------------------------------------------------
    localparam PKT_ADDR_H = 351;
    localparam PKT_ADDR_L = 288;
    localparam PKT_DEST_ID_H = 390;
    localparam PKT_DEST_ID_L = 386;
    localparam PKT_PROTECTION_H = 394;
    localparam PKT_PROTECTION_L = 392;
    localparam ST_DATA_W = 404;
    localparam ST_CHANNEL_W = 32;
    localparam DECODER_TYPE = 1;

    localparam PKT_TRANS_WRITE = 354;
    localparam PKT_TRANS_READ  = 355;

    localparam PKT_ADDR_W = PKT_ADDR_H-PKT_ADDR_L + 1;
    localparam PKT_DEST_ID_W = PKT_DEST_ID_H-PKT_DEST_ID_L + 1;



    // -------------------------------------------------------
    // Figure out the number of bits to mask off for each slave span
    // during address decoding
    // -------------------------------------------------------
    // -------------------------------------------------------
    // Work out which address bits are significant based on the
    // address range of the slaves. If the required width is too
    // large or too small, we use the address field width instead.
    // -------------------------------------------------------
    localparam ADDR_RANGE = 64'h0;
    localparam RANGE_ADDR_WIDTH = log2ceil(ADDR_RANGE);
    localparam OPTIMIZED_ADDR_H = (RANGE_ADDR_WIDTH > PKT_ADDR_W) ||
                                  (RANGE_ADDR_WIDTH == 0) ?
                                        PKT_ADDR_H :
                                        PKT_ADDR_L + RANGE_ADDR_WIDTH - 1;

    localparam RG = RANGE_ADDR_WIDTH;
    localparam REAL_ADDRESS_RANGE = OPTIMIZED_ADDR_H - PKT_ADDR_L;

    reg [PKT_DEST_ID_W-1 : 0] destid;

    // -------------------------------------------------------
    // Pass almost everything through, untouched
    // -------------------------------------------------------
    assign sink_ready        = src_ready;
    assign src_valid         = sink_valid;
    assign src_startofpacket = sink_startofpacket;
    assign src_endofpacket   = sink_endofpacket;
    wire [32-1 : 0] default_src_channel;




    // -------------------------------------------------------
    // Write and read transaction signals
    // -------------------------------------------------------
    wire read_transaction;
    assign read_transaction  = sink_data[PKT_TRANS_READ];


    MebX_Qsys_Project_mm_interconnect_0_router_032_default_decode the_default_decode(
      .default_destination_id (),
      .default_wr_channel   (),
      .default_rd_channel   (),
      .default_src_channel  (default_src_channel)
    );

    always @* begin
        src_data    = sink_data;
        src_channel = default_src_channel;

        // --------------------------------------------------
        // DestinationID Decoder
        // Sets the channel based on the destination ID.
        // --------------------------------------------------
        destid      = sink_data[PKT_DEST_ID_H : PKT_DEST_ID_L];



        if (destid == 24 ) begin
            src_channel = 32'b00000000000000000000000000000001;
        end

        if (destid == 0  && read_transaction) begin
            src_channel = 32'b00000000000000000000000000000010;
        end

        if (destid == 13 ) begin
            src_channel = 32'b00000000000000000000010000000000;
        end

        if (destid == 17 ) begin
            src_channel = 32'b00000000000000000000100000000000;
        end

        if (destid == 21 ) begin
            src_channel = 32'b00000000000000000001000000000000;
        end

        if (destid == 2  && read_transaction) begin
            src_channel = 32'b00000000000000000010000000000000;
        end

        if (destid == 6  && read_transaction) begin
            src_channel = 32'b00000000000000000100000000000000;
        end

        if (destid == 10  && read_transaction) begin
            src_channel = 32'b00000000000000001000000000000000;
        end

        if (destid == 14  && read_transaction) begin
            src_channel = 32'b00000000000000010000000000000000;
        end

        if (destid == 18  && read_transaction) begin
            src_channel = 32'b00000000000000100000000000000000;
        end

        if (destid == 22  && read_transaction) begin
            src_channel = 32'b00000000000001000000000000000000;
        end

        if (destid == 3 ) begin
            src_channel = 32'b00000000000010000000000000000000;
        end

        if (destid == 4  && read_transaction) begin
            src_channel = 32'b00000000000000000000000000000100;
        end

        if (destid == 7 ) begin
            src_channel = 32'b00000000000100000000000000000000;
        end

        if (destid == 11 ) begin
            src_channel = 32'b00000000001000000000000000000000;
        end

        if (destid == 15 ) begin
            src_channel = 32'b00000000010000000000000000000000;
        end

        if (destid == 23 ) begin
            src_channel = 32'b00000000100000000000000000000000;
        end

        if (destid == 19 ) begin
            src_channel = 32'b00000001000000000000000000000000;
        end

        if (destid == 26 ) begin
            src_channel = 32'b00000010000000000000000000000000;
        end

        if (destid == 27 ) begin
            src_channel = 32'b00000100000000000000000000000000;
        end

        if (destid == 28 ) begin
            src_channel = 32'b00001000000000000000000000000000;
        end

        if (destid == 29 ) begin
            src_channel = 32'b00010000000000000000000000000000;
        end

        if (destid == 30 ) begin
            src_channel = 32'b00100000000000000000000000000000;
        end

        if (destid == 8  && read_transaction) begin
            src_channel = 32'b00000000000000000000000000001000;
        end

        if (destid == 31 ) begin
            src_channel = 32'b01000000000000000000000000000000;
        end

        if (destid == 25 ) begin
            src_channel = 32'b10000000000000000000000000000000;
        end

        if (destid == 12  && read_transaction) begin
            src_channel = 32'b00000000000000000000000000010000;
        end

        if (destid == 16  && read_transaction) begin
            src_channel = 32'b00000000000000000000000000100000;
        end

        if (destid == 20  && read_transaction) begin
            src_channel = 32'b00000000000000000000000001000000;
        end

        if (destid == 1 ) begin
            src_channel = 32'b00000000000000000000000010000000;
        end

        if (destid == 5 ) begin
            src_channel = 32'b00000000000000000000000100000000;
        end

        if (destid == 9 ) begin
            src_channel = 32'b00000000000000000000001000000000;
        end


end


    // --------------------------------------------------
    // Ceil(log2()) function
    // --------------------------------------------------
    function integer log2ceil;
        input reg[65:0] val;
        reg [65:0] i;

        begin
            i = 1;
            log2ceil = 0;

            while (i < val) begin
                log2ceil = log2ceil + 1;
                i = i << 1;
            end
        end
    endfunction

endmodule


