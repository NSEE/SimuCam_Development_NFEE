io_out_5b_inst : io_out_5b PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig
	);
