spwr_select_in_altiobuf_inst : spwr_select_in_altiobuf PORT MAP (
		datain	 => datain_sig,
		dataout	 => dataout_sig
	);
