library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity comm_spw_mux_ent is
	port(
		-- basic inputs
		clk_i : in std_logic;
		rst_i : in std_logic
		-- logic inputs
		-- logic outputs
	);
end entity comm_spw_mux_ent;

architecture RTL of comm_spw_mux_ent is
	
begin

end architecture RTL;
