package comm_spw_codec_pkg is
	
end package comm_spw_codec_pkg;

package body comm_spw_codec_pkg is
	
end package body comm_spw_codec_pkg;
