library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity file is
	port(
		clk : in std_logic;
		rst : in std_logic
	);
end entity file;

architecture RTL of file is
	
begin

end architecture RTL;
