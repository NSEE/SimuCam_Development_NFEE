library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity testbench_top is
	port(
		clk : in std_logic;
		rst : in std_logic
	);
end entity testbench_top;

architecture RTL of testbench_top is
	
begin

end architecture RTL;
