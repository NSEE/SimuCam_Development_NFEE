library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity comm_v1_1_top is
	port(
		clk_i : in std_logic;
		rst_i : in std_logic
	);
end entity comm_v1_1_top;

architecture RTL of comm_v1_1_top is
	
	-- constants
	-- signals
	
begin
	
	-- spw codec instantiation
	
	-- spw mux/demux instantiation
	
	-- rmap codec instantiation
	
	-- rmap memory area instantiation
	
		
end architecture RTL;
